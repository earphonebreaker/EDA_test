
module dip_driver ( dip1, dip2, dip3, dip4, dip5, dip6, dip7, dip8, dip9, 
        reset_n, key1sel, key2sel, decrypt, desEnable, desIn );
  output [3:1] key1sel;
  output [3:1] key2sel;
  output [63:0] desIn;
  input dip1, dip2, dip3, dip4, dip5, dip6, dip7, dip8, dip9, reset_n;
  output decrypt, desEnable;
  wire   N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62,
         N63, N64, N65, N66, N67, N68, N71, N72, N73, N74, N75, N76, N77, N78,
         n2, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n3,
         n4, n5, n6, n7, n8, n9, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  OAI21X2 U13 ( .A0(n11), .A1(n12), .B0(n23), .Y(N68) );
  OAI21X2 U14 ( .A0(n12), .A1(n13), .B0(n23), .Y(N67) );
  OAI21X2 U15 ( .A0(n11), .A1(n14), .B0(n23), .Y(N66) );
  OAI21X2 U16 ( .A0(n13), .A1(n14), .B0(n23), .Y(N65) );
  OAI21X2 U17 ( .A0(n11), .A1(n15), .B0(n23), .Y(N64) );
  OAI21X2 U18 ( .A0(n13), .A1(n15), .B0(n23), .Y(N63) );
  OAI21X2 U19 ( .A0(n11), .A1(n16), .B0(n23), .Y(N62) );
  NAND2X2 U20 ( .A(n17), .B(dip5), .Y(n11) );
  OAI21X2 U21 ( .A0(n13), .A1(n16), .B0(n24), .Y(N61) );
  NAND2X2 U22 ( .A(n17), .B(n28), .Y(n13) );
  OAI21X2 U24 ( .A0(n12), .A1(n19), .B0(n24), .Y(N60) );
  OAI21X2 U25 ( .A0(n12), .A1(n20), .B0(n24), .Y(N59) );
  NAND2X2 U26 ( .A(dip6), .B(dip7), .Y(n12) );
  OAI21X2 U27 ( .A0(n14), .A1(n19), .B0(n24), .Y(N58) );
  OAI21X2 U28 ( .A0(n14), .A1(n20), .B0(n24), .Y(N57) );
  NAND2X2 U29 ( .A(dip7), .B(n29), .Y(n14) );
  OAI21X2 U30 ( .A0(n15), .A1(n19), .B0(n24), .Y(N56) );
  OAI21X2 U31 ( .A0(n15), .A1(n20), .B0(n24), .Y(N55) );
  NAND2X2 U32 ( .A(dip6), .B(n30), .Y(n15) );
  OAI21X2 U33 ( .A0(n16), .A1(n19), .B0(n24), .Y(N54) );
  NAND2X2 U34 ( .A(n21), .B(dip5), .Y(n19) );
  OAI21X2 U39 ( .A0(n16), .A1(n20), .B0(n23), .Y(N49) );
  NAND2X2 U40 ( .A(n21), .B(n28), .Y(n20) );
  NAND2X2 U43 ( .A(n29), .B(n30), .Y(n16) );
  TLATX1 \desIn_reg[63]  ( .G(N68), .D(n3), .Q(desIn[63]) );
  TLATX1 \desIn_reg[62]  ( .G(N68), .D(n4), .Q(desIn[62]) );
  TLATX1 \desIn_reg[61]  ( .G(N68), .D(n5), .Q(desIn[61]) );
  TLATX1 \desIn_reg[60]  ( .G(N68), .D(n6), .Q(desIn[60]) );
  TLATX1 \desIn_reg[59]  ( .G(N67), .D(n3), .Q(desIn[59]) );
  TLATX1 \desIn_reg[58]  ( .G(N67), .D(n4), .Q(desIn[58]) );
  TLATX1 \desIn_reg[57]  ( .G(N67), .D(n5), .Q(desIn[57]) );
  TLATX1 \desIn_reg[56]  ( .G(N67), .D(n6), .Q(desIn[56]) );
  TLATX1 \desIn_reg[55]  ( .G(N66), .D(n3), .Q(desIn[55]) );
  TLATX1 \desIn_reg[54]  ( .G(N66), .D(n4), .Q(desIn[54]) );
  TLATX1 \desIn_reg[53]  ( .G(N66), .D(n5), .Q(desIn[53]) );
  TLATX1 \desIn_reg[52]  ( .G(N66), .D(n6), .Q(desIn[52]) );
  TLATX1 \desIn_reg[51]  ( .G(N65), .D(n3), .Q(desIn[51]) );
  TLATX1 \desIn_reg[50]  ( .G(N65), .D(n4), .Q(desIn[50]) );
  TLATX1 \desIn_reg[49]  ( .G(N65), .D(n5), .Q(desIn[49]) );
  TLATX1 \desIn_reg[48]  ( .G(N65), .D(n6), .Q(desIn[48]) );
  TLATX1 \desIn_reg[47]  ( .G(N64), .D(n3), .Q(desIn[47]) );
  TLATX1 \desIn_reg[46]  ( .G(N64), .D(n4), .Q(desIn[46]) );
  TLATX1 \desIn_reg[45]  ( .G(N64), .D(n5), .Q(desIn[45]) );
  TLATX1 \desIn_reg[44]  ( .G(N64), .D(n6), .Q(desIn[44]) );
  TLATX1 \desIn_reg[43]  ( .G(N63), .D(n3), .Q(desIn[43]) );
  TLATX1 \desIn_reg[42]  ( .G(N63), .D(n4), .Q(desIn[42]) );
  TLATX1 \desIn_reg[41]  ( .G(N63), .D(n5), .Q(desIn[41]) );
  TLATX1 \desIn_reg[40]  ( .G(N63), .D(n6), .Q(desIn[40]) );
  TLATX1 \desIn_reg[39]  ( .G(N62), .D(n3), .Q(desIn[39]) );
  TLATX1 \desIn_reg[38]  ( .G(N62), .D(n4), .Q(desIn[38]) );
  TLATX1 \desIn_reg[37]  ( .G(N62), .D(n5), .Q(desIn[37]) );
  TLATX1 \desIn_reg[36]  ( .G(N62), .D(n6), .Q(desIn[36]) );
  TLATX1 \desIn_reg[35]  ( .G(N61), .D(n3), .Q(desIn[35]) );
  TLATX1 \desIn_reg[34]  ( .G(N61), .D(n4), .Q(desIn[34]) );
  TLATX1 \desIn_reg[33]  ( .G(N61), .D(n5), .Q(desIn[33]) );
  TLATX1 \desIn_reg[32]  ( .G(N61), .D(n6), .Q(desIn[32]) );
  TLATX1 \desIn_reg[31]  ( .G(N60), .D(n22), .Q(desIn[31]) );
  TLATX1 \desIn_reg[30]  ( .G(N60), .D(n9), .Q(desIn[30]) );
  TLATX1 \desIn_reg[29]  ( .G(N60), .D(n8), .Q(desIn[29]) );
  TLATX1 \desIn_reg[28]  ( .G(N60), .D(n7), .Q(desIn[28]) );
  TLATX1 \desIn_reg[27]  ( .G(N59), .D(n22), .Q(desIn[27]) );
  TLATX1 \desIn_reg[26]  ( .G(N59), .D(n9), .Q(desIn[26]) );
  TLATX1 \desIn_reg[25]  ( .G(N59), .D(n8), .Q(desIn[25]) );
  TLATX1 \desIn_reg[24]  ( .G(N59), .D(n7), .Q(desIn[24]) );
  TLATX1 \desIn_reg[23]  ( .G(N58), .D(n22), .Q(desIn[23]) );
  TLATX1 \desIn_reg[22]  ( .G(N58), .D(n9), .Q(desIn[22]) );
  TLATX1 \desIn_reg[21]  ( .G(N58), .D(n8), .Q(desIn[21]) );
  TLATX1 \desIn_reg[20]  ( .G(N58), .D(n7), .Q(desIn[20]) );
  TLATX1 \desIn_reg[19]  ( .G(N57), .D(n22), .Q(desIn[19]) );
  TLATX1 \desIn_reg[18]  ( .G(N57), .D(n9), .Q(desIn[18]) );
  TLATX1 \desIn_reg[17]  ( .G(N57), .D(n8), .Q(desIn[17]) );
  TLATX1 \desIn_reg[16]  ( .G(N57), .D(n7), .Q(desIn[16]) );
  TLATX1 \desIn_reg[15]  ( .G(N56), .D(n22), .Q(desIn[15]) );
  TLATX1 \desIn_reg[14]  ( .G(N56), .D(n9), .Q(desIn[14]) );
  TLATX1 \desIn_reg[13]  ( .G(N56), .D(n8), .Q(desIn[13]) );
  TLATX1 \desIn_reg[12]  ( .G(N56), .D(n7), .Q(desIn[12]) );
  TLATX1 \desIn_reg[11]  ( .G(N55), .D(n22), .Q(desIn[11]) );
  TLATX1 \desIn_reg[10]  ( .G(N55), .D(n9), .Q(desIn[10]) );
  TLATX1 \desIn_reg[9]  ( .G(N55), .D(n8), .Q(desIn[9]) );
  TLATX1 \desIn_reg[8]  ( .G(N55), .D(n7), .Q(desIn[8]) );
  TLATX1 \desIn_reg[7]  ( .G(N54), .D(n22), .Q(desIn[7]) );
  TLATX1 \desIn_reg[6]  ( .G(N54), .D(n9), .Q(desIn[6]) );
  TLATX1 \desIn_reg[5]  ( .G(N54), .D(n8), .Q(desIn[5]) );
  TLATX1 \desIn_reg[4]  ( .G(N54), .D(n7), .Q(desIn[4]) );
  TLATX1 \desIn_reg[3]  ( .G(N49), .D(n22), .Q(desIn[3]) );
  TLATX1 \desIn_reg[2]  ( .G(N49), .D(n9), .Q(desIn[2]) );
  TLATX1 \desIn_reg[1]  ( .G(N49), .D(n8), .Q(desIn[1]) );
  TLATX1 \desIn_reg[0]  ( .G(N49), .D(n7), .Q(desIn[0]) );
  TLATXL \key2sel_reg[3]  ( .G(N71), .D(N77), .Q(key2sel[3]) );
  TLATXL \key1sel_reg[3]  ( .G(N71), .D(N74), .Q(key1sel[3]) );
  TLATXL \key2sel_reg[2]  ( .G(N71), .D(N76), .Q(key2sel[2]) );
  TLATSRX1 desEnable_reg ( .G(dip9), .D(dip8), .RN(n23), .SN(1'b1), .Q(
        desEnable) );
  CLKINVX1 U44 ( .A(dip1), .Y(n2) );
  TLATXL decrypt_reg ( .G(N71), .D(N78), .Q(decrypt) );
  TLATXL \key1sel_reg[2]  ( .G(N71), .D(N73), .Q(key1sel[2]) );
  TLATXL \key2sel_reg[1]  ( .G(N71), .D(N75), .Q(key2sel[1]) );
  TLATXL \key1sel_reg[1]  ( .G(N71), .D(N72), .Q(key1sel[1]) );
  CLKBUFX4 U4 ( .A(reset_n), .Y(n23) );
  NAND2BX2 U5 ( .AN(dip9), .B(n23), .Y(n18) );
  CLKBUFX3 U6 ( .A(n22), .Y(n3) );
  CLKBUFX3 U7 ( .A(N53), .Y(n22) );
  CLKBUFX3 U8 ( .A(n9), .Y(n4) );
  CLKBUFX3 U9 ( .A(N52), .Y(n9) );
  CLKBUFX3 U10 ( .A(n8), .Y(n5) );
  CLKBUFX3 U11 ( .A(N51), .Y(n8) );
  CLKBUFX3 U12 ( .A(n7), .Y(n6) );
  CLKBUFX3 U23 ( .A(N50), .Y(n7) );
  OAI21X4 U35 ( .A0(dip8), .A1(n10), .B0(n24), .Y(N71) );
  NAND2X4 U36 ( .A(n24), .B(dip9), .Y(n10) );
  NOR2XL U37 ( .A(n10), .B(n2), .Y(N78) );
  NOR2XL U38 ( .A(n10), .B(n28), .Y(N75) );
  NOR2XL U41 ( .A(n10), .B(n29), .Y(N76) );
  NOR2XL U42 ( .A(n10), .B(n30), .Y(N77) );
  NOR2XL U45 ( .A(n10), .B(n25), .Y(N72) );
  NOR2XL U46 ( .A(n10), .B(n26), .Y(N73) );
  NOR2XL U47 ( .A(n10), .B(n27), .Y(N74) );
  NOR2X1 U48 ( .A(n2), .B(n18), .Y(N50) );
  NOR2X1 U49 ( .A(n25), .B(n18), .Y(N51) );
  NOR2X1 U50 ( .A(n26), .B(n18), .Y(N52) );
  NOR2X1 U51 ( .A(n27), .B(n18), .Y(N53) );
  NOR2X1 U52 ( .A(n18), .B(dip8), .Y(n21) );
  NOR2X1 U53 ( .A(n18), .B(n31), .Y(n17) );
  CLKINVX1 U54 ( .A(dip8), .Y(n31) );
  CLKINVX1 U55 ( .A(dip4), .Y(n27) );
  CLKINVX1 U56 ( .A(dip2), .Y(n25) );
  CLKINVX1 U57 ( .A(dip3), .Y(n26) );
  CLKINVX1 U58 ( .A(dip7), .Y(n30) );
  CLKINVX1 U59 ( .A(dip5), .Y(n28) );
  CLKINVX1 U60 ( .A(dip6), .Y(n29) );
  CLKBUFX6 U61 ( .A(reset_n), .Y(n24) );
endmodule


module keybox ( key1sel, key2sel, key1, key2 );
  input [2:0] key1sel;
  input [2:0] key2sel;
  output [55:0] key1;
  output [55:0] key2;
  wire   n3, n4;

  INVX1 U3 ( .A(1'b1), .Y(key2[0]) );
  INVX1 U5 ( .A(1'b1), .Y(key2[1]) );
  INVX1 U7 ( .A(1'b1), .Y(key2[2]) );
  INVX1 U9 ( .A(1'b1), .Y(key2[3]) );
  INVX1 U11 ( .A(1'b1), .Y(key2[4]) );
  INVX1 U13 ( .A(1'b1), .Y(key2[5]) );
  INVX1 U15 ( .A(1'b1), .Y(key2[6]) );
  INVX1 U17 ( .A(1'b1), .Y(key2[7]) );
  INVX1 U19 ( .A(1'b1), .Y(key2[8]) );
  INVX1 U21 ( .A(1'b1), .Y(key2[9]) );
  INVX1 U23 ( .A(1'b1), .Y(key2[10]) );
  INVX1 U25 ( .A(1'b1), .Y(key2[11]) );
  INVX1 U27 ( .A(1'b1), .Y(key2[12]) );
  INVX1 U29 ( .A(1'b1), .Y(key2[13]) );
  INVX1 U31 ( .A(1'b1), .Y(key2[14]) );
  INVX1 U33 ( .A(1'b1), .Y(key2[15]) );
  INVX1 U35 ( .A(1'b1), .Y(key2[16]) );
  INVX1 U37 ( .A(1'b1), .Y(key2[17]) );
  INVX1 U39 ( .A(1'b1), .Y(key2[18]) );
  INVX1 U41 ( .A(1'b1), .Y(key2[19]) );
  INVX1 U43 ( .A(1'b1), .Y(key2[20]) );
  INVX1 U45 ( .A(1'b1), .Y(key2[21]) );
  INVX1 U47 ( .A(1'b1), .Y(key2[22]) );
  INVX1 U49 ( .A(1'b1), .Y(key2[23]) );
  INVX1 U51 ( .A(1'b1), .Y(key2[24]) );
  INVX1 U53 ( .A(1'b1), .Y(key2[25]) );
  INVX1 U55 ( .A(1'b1), .Y(key2[26]) );
  INVX1 U57 ( .A(1'b1), .Y(key2[27]) );
  INVX1 U59 ( .A(1'b1), .Y(key2[28]) );
  INVX1 U61 ( .A(1'b1), .Y(key2[29]) );
  INVX1 U63 ( .A(1'b1), .Y(key2[30]) );
  INVX1 U65 ( .A(1'b1), .Y(key2[31]) );
  INVX1 U67 ( .A(1'b1), .Y(key2[32]) );
  INVX1 U69 ( .A(1'b1), .Y(key2[33]) );
  INVX1 U71 ( .A(1'b1), .Y(key2[34]) );
  INVX1 U73 ( .A(1'b1), .Y(key2[35]) );
  INVX1 U75 ( .A(1'b1), .Y(key2[36]) );
  INVX1 U77 ( .A(1'b1), .Y(key2[37]) );
  INVX1 U79 ( .A(1'b1), .Y(key2[38]) );
  INVX1 U81 ( .A(1'b1), .Y(key2[39]) );
  INVX1 U83 ( .A(1'b1), .Y(key2[40]) );
  INVX1 U85 ( .A(1'b1), .Y(key2[41]) );
  INVX1 U87 ( .A(1'b1), .Y(key2[42]) );
  INVX1 U89 ( .A(1'b1), .Y(key2[43]) );
  INVX1 U91 ( .A(1'b1), .Y(key2[48]) );
  INVX1 U93 ( .A(1'b1), .Y(key2[49]) );
  INVX1 U95 ( .A(1'b1), .Y(key2[50]) );
  INVX1 U97 ( .A(1'b1), .Y(key2[51]) );
  INVX1 U99 ( .A(1'b1), .Y(key2[52]) );
  INVX1 U101 ( .A(1'b1), .Y(key2[53]) );
  INVX1 U103 ( .A(1'b1), .Y(key2[54]) );
  INVX1 U105 ( .A(1'b1), .Y(key2[55]) );
  INVX1 U107 ( .A(1'b1), .Y(key1[0]) );
  INVX1 U109 ( .A(1'b1), .Y(key1[1]) );
  INVX1 U111 ( .A(1'b1), .Y(key1[2]) );
  INVX1 U113 ( .A(1'b1), .Y(key1[3]) );
  INVX1 U115 ( .A(1'b1), .Y(key1[4]) );
  INVX1 U117 ( .A(1'b1), .Y(key1[5]) );
  INVX1 U119 ( .A(1'b1), .Y(key1[6]) );
  INVX1 U121 ( .A(1'b1), .Y(key1[7]) );
  INVX1 U123 ( .A(1'b1), .Y(key1[8]) );
  INVX1 U125 ( .A(1'b1), .Y(key1[9]) );
  INVX1 U127 ( .A(1'b1), .Y(key1[10]) );
  INVX1 U129 ( .A(1'b1), .Y(key1[11]) );
  INVX1 U131 ( .A(1'b1), .Y(key1[12]) );
  INVX1 U133 ( .A(1'b1), .Y(key1[13]) );
  INVX1 U135 ( .A(1'b1), .Y(key1[14]) );
  INVX1 U137 ( .A(1'b1), .Y(key1[15]) );
  INVX1 U139 ( .A(1'b1), .Y(key1[16]) );
  INVX1 U141 ( .A(1'b1), .Y(key1[17]) );
  INVX1 U143 ( .A(1'b1), .Y(key1[18]) );
  INVX1 U145 ( .A(1'b1), .Y(key1[19]) );
  INVX1 U147 ( .A(1'b1), .Y(key1[20]) );
  INVX1 U149 ( .A(1'b1), .Y(key1[21]) );
  INVX1 U151 ( .A(1'b1), .Y(key1[22]) );
  INVX1 U153 ( .A(1'b1), .Y(key1[23]) );
  INVX1 U155 ( .A(1'b1), .Y(key1[24]) );
  INVX1 U157 ( .A(1'b1), .Y(key1[25]) );
  INVX1 U159 ( .A(1'b1), .Y(key1[26]) );
  INVX1 U161 ( .A(1'b1), .Y(key1[27]) );
  INVX1 U163 ( .A(1'b1), .Y(key1[28]) );
  INVX1 U165 ( .A(1'b1), .Y(key1[29]) );
  INVX1 U167 ( .A(1'b1), .Y(key1[30]) );
  INVX1 U169 ( .A(1'b1), .Y(key1[31]) );
  INVX1 U171 ( .A(1'b1), .Y(key1[32]) );
  INVX1 U173 ( .A(1'b1), .Y(key1[33]) );
  INVX1 U175 ( .A(1'b1), .Y(key1[34]) );
  INVX1 U177 ( .A(1'b1), .Y(key1[35]) );
  INVX1 U179 ( .A(1'b1), .Y(key1[36]) );
  INVX1 U181 ( .A(1'b1), .Y(key1[37]) );
  INVX1 U183 ( .A(1'b1), .Y(key1[38]) );
  INVX1 U185 ( .A(1'b1), .Y(key1[39]) );
  INVX1 U187 ( .A(1'b1), .Y(key1[40]) );
  INVX1 U189 ( .A(1'b1), .Y(key1[41]) );
  INVX1 U191 ( .A(1'b1), .Y(key1[42]) );
  INVX1 U193 ( .A(1'b1), .Y(key1[43]) );
  INVX1 U195 ( .A(1'b1), .Y(key1[48]) );
  INVX1 U197 ( .A(1'b1), .Y(key1[49]) );
  INVX1 U199 ( .A(1'b1), .Y(key1[50]) );
  INVX1 U201 ( .A(1'b1), .Y(key1[51]) );
  INVX1 U203 ( .A(1'b1), .Y(key1[52]) );
  INVX1 U205 ( .A(1'b1), .Y(key1[53]) );
  INVX1 U207 ( .A(1'b1), .Y(key1[54]) );
  INVX1 U209 ( .A(1'b1), .Y(key1[55]) );
  NAND2X1 U211 ( .A(key2sel[1]), .B(key2sel[0]), .Y(n3) );
  NAND2X1 U212 ( .A(key1sel[1]), .B(key1sel[0]), .Y(n4) );
  CLKINVX1 U213 ( .A(key2sel[0]), .Y(key2[44]) );
  CLKINVX1 U214 ( .A(key1sel[0]), .Y(key1[44]) );
  XOR2X1 U215 ( .A(key2sel[1]), .B(key2sel[0]), .Y(key2[45]) );
  XOR2X1 U216 ( .A(key1sel[1]), .B(key1sel[0]), .Y(key1[45]) );
  XNOR2X1 U217 ( .A(key2sel[2]), .B(n3), .Y(key2[46]) );
  XNOR2X1 U218 ( .A(key1sel[2]), .B(n4), .Y(key1[46]) );
  AND3X2 U219 ( .A(key1sel[2]), .B(key1sel[0]), .C(key1sel[1]), .Y(key1[47])
         );
  NOR2BX1 U220 ( .AN(key2sel[2]), .B(n3), .Y(key2[47]) );
endmodule


module key_sel ( clk, K, decrypt, K1, K2, K3, K4, K5, K6, K7, K8, K9, K10, K11, 
        K12, K13, K14, K15, K16 );
  input [55:0] K;
  output [1:48] K1;
  output [1:48] K2;
  output [1:48] K3;
  output [1:48] K4;
  output [1:48] K5;
  output [1:48] K6;
  output [1:48] K7;
  output [1:48] K8;
  output [1:48] K9;
  output [1:48] K10;
  output [1:48] K11;
  output [1:48] K12;
  output [1:48] K13;
  output [1:48] K14;
  output [1:48] K15;
  output [1:48] K16;
  input clk, decrypt;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433;
  wire   [55:0] K_r0;
  wire   [55:0] K_r1;
  wire   [55:0] K_r2;
  wire   [55:0] K_r3;
  wire   [55:0] K_r4;
  wire   [55:0] K_r5;
  wire   [55:0] K_r6;
  wire   [55:0] K_r7;
  wire   [55:0] K_r8;
  wire   [55:0] K_r9;
  wire   [55:0] K_r10;
  wire   [55:0] K_r11;
  wire   [55:0] K_r12;
  wire   [55:0] K_r14;
  wire   [55:0] K_r13;

  DFFQX1 \K_r14_reg[50]  ( .D(K_r13[50]), .CK(n278), .Q(K_r14[50]) );
  DFFQX1 \K_r14_reg[49]  ( .D(K_r13[49]), .CK(n278), .Q(K_r14[49]) );
  DFFQX1 \K_r14_reg[46]  ( .D(K_r13[46]), .CK(n278), .Q(K_r14[46]) );
  DFFQX1 \K_r14_reg[45]  ( .D(K_r13[45]), .CK(n278), .Q(K_r14[45]) );
  DFFQX1 \K_r14_reg[43]  ( .D(K_r13[43]), .CK(n277), .Q(K_r14[43]) );
  DFFQX1 \K_r14_reg[42]  ( .D(K_r13[42]), .CK(n277), .Q(K_r14[42]) );
  DFFQX1 \K_r14_reg[39]  ( .D(K_r13[39]), .CK(n277), .Q(K_r14[39]) );
  DFFQX1 \K_r14_reg[38]  ( .D(K_r13[38]), .CK(n277), .Q(K_r14[38]) );
  DFFQX1 \K_r14_reg[18]  ( .D(K_r13[18]), .CK(n275), .Q(K_r14[18]) );
  DFFQX1 \K_r14_reg[15]  ( .D(K_r13[15]), .CK(n274), .Q(K_r14[15]) );
  DFFQX1 \K_r14_reg[12]  ( .D(K_r13[12]), .CK(n274), .Q(K_r14[12]) );
  DFFQX1 \K_r14_reg[11]  ( .D(K_r13[11]), .CK(n274), .Q(K_r14[11]) );
  DFFQX1 \K_r14_reg[10]  ( .D(K_r13[10]), .CK(n274), .Q(K_r14[10]) );
  DFFQX1 \K_r14_reg[8]  ( .D(K_r13[8]), .CK(n273), .Q(K_r14[8]) );
  DFFQX1 \K_r14_reg[5]  ( .D(K_r13[5]), .CK(n273), .Q(K_r14[5]) );
  DFFQX1 \K_r14_reg[3]  ( .D(K_r13[3]), .CK(n273), .Q(K_r14[3]) );
  DFFQX1 \K_r6_reg[55]  ( .D(K_r5[55]), .CK(n340), .Q(K_r6[55]) );
  DFFQX1 \K_r7_reg[55]  ( .D(K_r6[55]), .CK(n340), .Q(K_r7[55]) );
  DFFQX1 \K_r13_reg[55]  ( .D(K_r12[55]), .CK(n339), .Q(K_r13[55]) );
  DFFQX1 \K_r4_reg[54]  ( .D(K_r3[54]), .CK(n339), .Q(K_r4[54]) );
  DFFQX1 \K_r9_reg[54]  ( .D(K_r8[54]), .CK(n338), .Q(K_r9[54]) );
  DFFQX1 \K_r2_reg[53]  ( .D(K_r1[53]), .CK(n337), .Q(K_r2[53]) );
  DFFQX1 \K_r6_reg[53]  ( .D(K_r5[53]), .CK(n337), .Q(K_r6[53]) );
  DFFQX1 \K_r7_reg[53]  ( .D(K_r6[53]), .CK(n337), .Q(K_r7[53]) );
  DFFQX1 \K_r11_reg[53]  ( .D(K_r10[53]), .CK(n336), .Q(K_r11[53]) );
  DFFQX1 \K_r0_reg[52]  ( .D(K[52]), .CK(n336), .Q(K_r0[52]) );
  DFFQX1 \K_r3_reg[52]  ( .D(K_r2[52]), .CK(n336), .Q(K_r3[52]) );
  DFFQX1 \K_r10_reg[52]  ( .D(K_r9[52]), .CK(n335), .Q(K_r10[52]) );
  DFFQX1 \K_r13_reg[52]  ( .D(K_r12[52]), .CK(n335), .Q(K_r13[52]) );
  DFFQX1 \K_r5_reg[51]  ( .D(K_r4[51]), .CK(n334), .Q(K_r5[51]) );
  DFFQX1 \K_r6_reg[51]  ( .D(K_r5[51]), .CK(n334), .Q(K_r6[51]) );
  DFFQX1 \K_r7_reg[51]  ( .D(K_r6[51]), .CK(n334), .Q(K_r7[51]) );
  DFFQX1 \K_r8_reg[51]  ( .D(K_r7[51]), .CK(n334), .Q(K_r8[51]) );
  DFFQX1 \K_r2_reg[50]  ( .D(K_r1[50]), .CK(n333), .Q(K_r2[50]) );
  DFFQX1 \K_r11_reg[50]  ( .D(K_r10[50]), .CK(n332), .Q(K_r11[50]) );
  DFFQX1 \K_r3_reg[49]  ( .D(K_r2[49]), .CK(n331), .Q(K_r3[49]) );
  DFFQX1 \K_r4_reg[49]  ( .D(K_r3[49]), .CK(n331), .Q(K_r4[49]) );
  DFFQX1 \K_r9_reg[49]  ( .D(K_r8[49]), .CK(n330), .Q(K_r9[49]) );
  DFFQX1 \K_r10_reg[49]  ( .D(K_r9[49]), .CK(n330), .Q(K_r10[49]) );
  DFFQX1 \K_r4_reg[48]  ( .D(K_r3[48]), .CK(n329), .Q(K_r4[48]) );
  DFFQX1 \K_r5_reg[48]  ( .D(K_r4[48]), .CK(n329), .Q(K_r5[48]) );
  DFFQX1 \K_r8_reg[48]  ( .D(K_r7[48]), .CK(n329), .Q(K_r8[48]) );
  DFFQX1 \K_r9_reg[48]  ( .D(K_r8[48]), .CK(n329), .Q(K_r9[48]) );
  DFFQX1 \K_r1_reg[47]  ( .D(K_r0[47]), .CK(n328), .Q(K_r1[47]) );
  DFFQX1 \K_r2_reg[47]  ( .D(K_r1[47]), .CK(n328), .Q(K_r2[47]) );
  DFFQX1 \K_r3_reg[47]  ( .D(K_r2[47]), .CK(n328), .Q(K_r3[47]) );
  DFFQX1 \K_r10_reg[47]  ( .D(K_r9[47]), .CK(n327), .Q(K_r10[47]) );
  DFFQX1 \K_r11_reg[47]  ( .D(K_r10[47]), .CK(n327), .Q(K_r11[47]) );
  DFFQX1 \K_r12_reg[47]  ( .D(K_r11[47]), .CK(n327), .Q(K_r12[47]) );
  DFFQX1 \K_r6_reg[46]  ( .D(K_r5[46]), .CK(n326), .Q(K_r6[46]) );
  DFFQX1 \K_r7_reg[46]  ( .D(K_r6[46]), .CK(n326), .Q(K_r7[46]) );
  DFFQX1 \K_r1_reg[44]  ( .D(K_r0[44]), .CK(n324), .Q(K_r1[44]) );
  DFFQX1 \K_r3_reg[44]  ( .D(K_r2[44]), .CK(n323), .Q(K_r3[44]) );
  DFFQX1 \K_r10_reg[44]  ( .D(K_r9[44]), .CK(n323), .Q(K_r10[44]) );
  DFFQX1 \K_r12_reg[44]  ( .D(K_r11[44]), .CK(n322), .Q(K_r12[44]) );
  DFFQX1 \K_r3_reg[43]  ( .D(K_r2[43]), .CK(n322), .Q(K_r3[43]) );
  DFFQX1 \K_r5_reg[43]  ( .D(K_r4[43]), .CK(n322), .Q(K_r5[43]) );
  DFFQX1 \K_r8_reg[43]  ( .D(K_r7[43]), .CK(n321), .Q(K_r8[43]) );
  DFFQX1 \K_r10_reg[43]  ( .D(K_r9[43]), .CK(n321), .Q(K_r10[43]) );
  DFFQX1 \K_r1_reg[42]  ( .D(K_r0[42]), .CK(n320), .Q(K_r1[42]) );
  DFFQX1 \K_r12_reg[42]  ( .D(K_r11[42]), .CK(n319), .Q(K_r12[42]) );
  DFFQX1 \K_r1_reg[41]  ( .D(K_r0[41]), .CK(n319), .Q(K_r1[41]) );
  DFFQX1 \K_r5_reg[41]  ( .D(K_r4[41]), .CK(n318), .Q(K_r5[41]) );
  DFFQX1 \K_r8_reg[41]  ( .D(K_r7[41]), .CK(n318), .Q(K_r8[41]) );
  DFFQX1 \K_r12_reg[41]  ( .D(K_r11[41]), .CK(n318), .Q(K_r12[41]) );
  DFFQX1 \K_r5_reg[40]  ( .D(K_r4[40]), .CK(n317), .Q(K_r5[40]) );
  DFFQX1 \K_r8_reg[40]  ( .D(K_r7[40]), .CK(n317), .Q(K_r8[40]) );
  DFFQX1 \K_r4_reg[38]  ( .D(K_r3[38]), .CK(n314), .Q(K_r4[38]) );
  DFFQX1 \K_r9_reg[38]  ( .D(K_r8[38]), .CK(n313), .Q(K_r9[38]) );
  DFFQX1 \K_r5_reg[37]  ( .D(K_r4[37]), .CK(n312), .Q(K_r5[37]) );
  DFFQX1 \K_r6_reg[37]  ( .D(K_r5[37]), .CK(n312), .Q(K_r6[37]) );
  DFFQX1 \K_r7_reg[37]  ( .D(K_r6[37]), .CK(n312), .Q(K_r7[37]) );
  DFFQX1 \K_r8_reg[37]  ( .D(K_r7[37]), .CK(n312), .Q(K_r8[37]) );
  DFFQX1 \K_r0_reg[36]  ( .D(K[36]), .CK(n311), .Q(K_r0[36]) );
  DFFQX1 \K_r1_reg[36]  ( .D(K_r0[36]), .CK(n311), .Q(K_r1[36]) );
  DFFQX1 \K_r12_reg[36]  ( .D(K_r11[36]), .CK(n310), .Q(K_r12[36]) );
  DFFQX1 \K_r13_reg[36]  ( .D(K_r12[36]), .CK(n310), .Q(K_r13[36]) );
  DFFQX1 \K_r0_reg[35]  ( .D(K[35]), .CK(n310), .Q(K_r0[35]) );
  DFFQX1 \K_r3_reg[35]  ( .D(K_r2[35]), .CK(n309), .Q(K_r3[35]) );
  DFFQX1 \K_r4_reg[35]  ( .D(K_r3[35]), .CK(n309), .Q(K_r4[35]) );
  DFFQX1 \K_r9_reg[35]  ( .D(K_r8[35]), .CK(n309), .Q(K_r9[35]) );
  DFFQX1 \K_r10_reg[35]  ( .D(K_r9[35]), .CK(n309), .Q(K_r10[35]) );
  DFFQX1 \K_r13_reg[35]  ( .D(K_r12[35]), .CK(n308), .Q(K_r13[35]) );
  DFFQX1 \K_r3_reg[34]  ( .D(K_r2[34]), .CK(n308), .Q(K_r3[34]) );
  DFFQX1 \K_r6_reg[34]  ( .D(K_r5[34]), .CK(n307), .Q(K_r6[34]) );
  DFFQX1 \K_r7_reg[34]  ( .D(K_r6[34]), .CK(n307), .Q(K_r7[34]) );
  DFFQX1 \K_r10_reg[34]  ( .D(K_r9[34]), .CK(n307), .Q(K_r10[34]) );
  DFFQX1 \K_r1_reg[33]  ( .D(K_r0[33]), .CK(n306), .Q(K_r1[33]) );
  DFFQX1 \K_r2_reg[33]  ( .D(K_r1[33]), .CK(n306), .Q(K_r2[33]) );
  DFFQX1 \K_r4_reg[33]  ( .D(K_r3[33]), .CK(n306), .Q(K_r4[33]) );
  DFFQX1 \K_r9_reg[33]  ( .D(K_r8[33]), .CK(n306), .Q(K_r9[33]) );
  DFFQX1 \K_r11_reg[33]  ( .D(K_r10[33]), .CK(n305), .Q(K_r11[33]) );
  DFFQX1 \K_r12_reg[33]  ( .D(K_r11[33]), .CK(n305), .Q(K_r12[33]) );
  DFFQX1 \K_r0_reg[32]  ( .D(K[32]), .CK(n305), .Q(K_r0[32]) );
  DFFQX1 \K_r5_reg[32]  ( .D(K_r4[32]), .CK(n304), .Q(K_r5[32]) );
  DFFQX1 \K_r8_reg[32]  ( .D(K_r7[32]), .CK(n304), .Q(K_r8[32]) );
  DFFQX1 \K_r13_reg[32]  ( .D(K_r12[32]), .CK(n304), .Q(K_r13[32]) );
  DFFQX1 \K_r0_reg[31]  ( .D(K[31]), .CK(n303), .Q(K_r0[31]) );
  DFFQX1 \K_r4_reg[31]  ( .D(K_r3[31]), .CK(n303), .Q(K_r4[31]) );
  DFFQX1 \K_r6_reg[31]  ( .D(K_r5[31]), .CK(n303), .Q(K_r6[31]) );
  DFFQX1 \K_r7_reg[31]  ( .D(K_r6[31]), .CK(n303), .Q(K_r7[31]) );
  DFFQX1 \K_r9_reg[31]  ( .D(K_r8[31]), .CK(n302), .Q(K_r9[31]) );
  DFFQX1 \K_r13_reg[31]  ( .D(K_r12[31]), .CK(n302), .Q(K_r13[31]) );
  DFFQX1 \K_r6_reg[30]  ( .D(K_r5[30]), .CK(n301), .Q(K_r6[30]) );
  DFFQX1 \K_r7_reg[30]  ( .D(K_r6[30]), .CK(n301), .Q(K_r7[30]) );
  DFFQX1 \K_r2_reg[29]  ( .D(K_r1[29]), .CK(n300), .Q(K_r2[29]) );
  DFFQX1 \K_r6_reg[29]  ( .D(K_r5[29]), .CK(n300), .Q(K_r6[29]) );
  DFFQX1 \K_r7_reg[29]  ( .D(K_r6[29]), .CK(n300), .Q(K_r7[29]) );
  DFFQX1 \K_r11_reg[29]  ( .D(K_r10[29]), .CK(n299), .Q(K_r11[29]) );
  DFFQX1 \K_r2_reg[28]  ( .D(K_r1[28]), .CK(n299), .Q(K_r2[28]) );
  DFFQX1 \K_r11_reg[28]  ( .D(K_r10[28]), .CK(n298), .Q(K_r11[28]) );
  DFFQX1 \K_r2_reg[27]  ( .D(K_r1[27]), .CK(n297), .Q(K_r2[27]) );
  DFFQX1 \K_r4_reg[27]  ( .D(K_r3[27]), .CK(n297), .Q(K_r4[27]) );
  DFFQX1 \K_r6_reg[27]  ( .D(K_r5[27]), .CK(n297), .Q(K_r6[27]) );
  DFFQX1 \K_r7_reg[27]  ( .D(K_r6[27]), .CK(n296), .Q(K_r7[27]) );
  DFFQX1 \K_r9_reg[27]  ( .D(K_r8[27]), .CK(n296), .Q(K_r9[27]) );
  DFFQX1 \K_r11_reg[27]  ( .D(K_r10[27]), .CK(n296), .Q(K_r11[27]) );
  DFFQX1 \K_r6_reg[26]  ( .D(K_r5[26]), .CK(n295), .Q(K_r6[26]) );
  DFFQX1 \K_r7_reg[26]  ( .D(K_r6[26]), .CK(n295), .Q(K_r7[26]) );
  DFFQX1 \K_r0_reg[25]  ( .D(K[25]), .CK(n294), .Q(K_r0[25]) );
  DFFQX1 \K_r2_reg[25]  ( .D(K_r1[25]), .CK(n294), .Q(K_r2[25]) );
  DFFQX1 \K_r11_reg[25]  ( .D(K_r10[25]), .CK(n293), .Q(K_r11[25]) );
  DFFQX1 \K_r13_reg[25]  ( .D(K_r12[25]), .CK(n293), .Q(K_r13[25]) );
  DFFQX1 \K_r2_reg[24]  ( .D(K_r1[24]), .CK(n292), .Q(K_r2[24]) );
  DFFQX1 \K_r11_reg[24]  ( .D(K_r10[24]), .CK(n291), .Q(K_r11[24]) );
  DFFQX1 \K_r4_reg[23]  ( .D(K_r3[23]), .CK(n291), .Q(K_r4[23]) );
  DFFQX1 \K_r9_reg[23]  ( .D(K_r8[23]), .CK(n290), .Q(K_r9[23]) );
  DFFQX1 \K_r0_reg[22]  ( .D(K[22]), .CK(n289), .Q(K_r0[22]) );
  DFFQX1 \K_r1_reg[22]  ( .D(K_r0[22]), .CK(n289), .Q(K_r1[22]) );
  DFFQX1 \K_r6_reg[22]  ( .D(K_r5[22]), .CK(n289), .Q(K_r6[22]) );
  DFFQX1 \K_r7_reg[22]  ( .D(K_r6[22]), .CK(n289), .Q(K_r7[22]) );
  DFFQX1 \K_r12_reg[22]  ( .D(K_r11[22]), .CK(n288), .Q(K_r12[22]) );
  DFFQX1 \K_r13_reg[22]  ( .D(K_r12[22]), .CK(n288), .Q(K_r13[22]) );
  DFFQX1 \K_r1_reg[21]  ( .D(K_r0[21]), .CK(n288), .Q(K_r1[21]) );
  DFFQX1 \K_r2_reg[21]  ( .D(K_r1[21]), .CK(n288), .Q(K_r2[21]) );
  DFFQX1 \K_r5_reg[21]  ( .D(K_r4[21]), .CK(n287), .Q(K_r5[21]) );
  DFFQX1 \K_r8_reg[21]  ( .D(K_r7[21]), .CK(n287), .Q(K_r8[21]) );
  DFFQX1 \K_r11_reg[21]  ( .D(K_r10[21]), .CK(n287), .Q(K_r11[21]) );
  DFFQX1 \K_r12_reg[21]  ( .D(K_r11[21]), .CK(n287), .Q(K_r12[21]) );
  DFFQX1 \K_r2_reg[20]  ( .D(K_r1[20]), .CK(n286), .Q(K_r2[20]) );
  DFFQX1 \K_r11_reg[20]  ( .D(K_r10[20]), .CK(n285), .Q(K_r11[20]) );
  DFFQX1 \K_r0_reg[19]  ( .D(K[19]), .CK(n285), .Q(K_r0[19]) );
  DFFQX1 \K_r3_reg[19]  ( .D(K_r2[19]), .CK(n284), .Q(K_r3[19]) );
  DFFQX1 \K_r5_reg[19]  ( .D(K_r4[19]), .CK(n284), .Q(K_r5[19]) );
  DFFQX1 \K_r6_reg[19]  ( .D(K_r5[19]), .CK(n284), .Q(K_r6[19]) );
  DFFQX1 \K_r7_reg[19]  ( .D(K_r6[19]), .CK(n284), .Q(K_r7[19]) );
  DFFQX1 \K_r8_reg[19]  ( .D(K_r7[19]), .CK(n284), .Q(K_r8[19]) );
  DFFQX1 \K_r10_reg[19]  ( .D(K_r9[19]), .CK(n284), .Q(K_r10[19]) );
  DFFQX1 \K_r13_reg[19]  ( .D(K_r12[19]), .CK(n283), .Q(K_r13[19]) );
  DFFQX1 \K_r1_reg[18]  ( .D(K_r0[18]), .CK(n283), .Q(K_r1[18]) );
  DFFQX1 \K_r4_reg[18]  ( .D(K_r3[18]), .CK(n283), .Q(K_r4[18]) );
  DFFQX1 \K_r9_reg[18]  ( .D(K_r8[18]), .CK(n282), .Q(K_r9[18]) );
  DFFQX1 \K_r12_reg[18]  ( .D(K_r11[18]), .CK(n282), .Q(K_r12[18]) );
  DFFQX1 \K_r0_reg[17]  ( .D(K[17]), .CK(n282), .Q(K_r0[17]) );
  DFFQX1 \K_r13_reg[17]  ( .D(K_r12[17]), .CK(n280), .Q(K_r13[17]) );
  DFFQX1 \K_r1_reg[16]  ( .D(K_r0[16]), .CK(n280), .Q(K_r1[16]) );
  DFFQX1 \K_r3_reg[16]  ( .D(K_r2[16]), .CK(n280), .Q(K_r3[16]) );
  DFFQX1 \K_r5_reg[16]  ( .D(K_r4[16]), .CK(n280), .Q(K_r5[16]) );
  DFFQX1 \K_r8_reg[16]  ( .D(K_r7[16]), .CK(n372), .Q(K_r8[16]) );
  DFFQX1 \K_r10_reg[16]  ( .D(K_r9[16]), .CK(n341), .Q(K_r10[16]) );
  DFFQX1 \K_r12_reg[16]  ( .D(K_r11[16]), .CK(n364), .Q(K_r12[16]) );
  DFFQX1 \K_r1_reg[15]  ( .D(K_r0[15]), .CK(n354), .Q(K_r1[15]) );
  DFFQX1 \K_r12_reg[15]  ( .D(K_r11[15]), .CK(n348), .Q(K_r12[15]) );
  DFFQX1 \K_r3_reg[14]  ( .D(K_r2[14]), .CK(n349), .Q(K_r3[14]) );
  DFFQX1 \K_r10_reg[14]  ( .D(K_r9[14]), .CK(n361), .Q(K_r10[14]) );
  DFFQX1 \K_r5_reg[13]  ( .D(K_r4[13]), .CK(n354), .Q(K_r5[13]) );
  DFFQX1 \K_r8_reg[13]  ( .D(K_r7[13]), .CK(n355), .Q(K_r8[13]) );
  DFFQX1 \K_r3_reg[11]  ( .D(K_r2[11]), .CK(n353), .Q(K_r3[11]) );
  DFFQX1 \K_r10_reg[11]  ( .D(K_r9[11]), .CK(n347), .Q(K_r10[11]) );
  DFFQX1 \K_r1_reg[10]  ( .D(K_r0[10]), .CK(n348), .Q(K_r1[10]) );
  DFFQX1 \K_r3_reg[10]  ( .D(K_r2[10]), .CK(n360), .Q(K_r3[10]) );
  DFFQX1 \K_r5_reg[10]  ( .D(K_r4[10]), .CK(n361), .Q(K_r5[10]) );
  DFFQX1 \K_r8_reg[10]  ( .D(K_r7[10]), .CK(n366), .Q(K_r8[10]) );
  DFFQX1 \K_r10_reg[10]  ( .D(K_r9[10]), .CK(n343), .Q(K_r10[10]) );
  DFFQX1 \K_r12_reg[10]  ( .D(K_r11[10]), .CK(n358), .Q(K_r12[10]) );
  DFFQX1 \K_r3_reg[9]  ( .D(K_r2[9]), .CK(n367), .Q(K_r3[9]) );
  DFFQX1 \K_r10_reg[9]  ( .D(K_r9[9]), .CK(n351), .Q(K_r10[9]) );
  DFFQX1 \K_r2_reg[8]  ( .D(K_r1[8]), .CK(n344), .Q(K_r2[8]) );
  DFFQX1 \K_r5_reg[8]  ( .D(K_r4[8]), .CK(n345), .Q(K_r5[8]) );
  DFFQX1 \K_r8_reg[8]  ( .D(K_r7[8]), .CK(n346), .Q(K_r8[8]) );
  DFFQX1 \K_r11_reg[8]  ( .D(K_r10[8]), .CK(n361), .Q(K_r11[8]) );
  DFFQX1 \K_r1_reg[7]  ( .D(K_r0[7]), .CK(n366), .Q(K_r1[7]) );
  DFFQX1 \K_r2_reg[7]  ( .D(K_r1[7]), .CK(n365), .Q(K_r2[7]) );
  DFFQX1 \K_r6_reg[7]  ( .D(K_r5[7]), .CK(n365), .Q(K_r6[7]) );
  DFFQX1 \K_r7_reg[7]  ( .D(K_r6[7]), .CK(n364), .Q(K_r7[7]) );
  DFFQX1 \K_r11_reg[7]  ( .D(K_r10[7]), .CK(n372), .Q(K_r11[7]) );
  DFFQX1 \K_r12_reg[7]  ( .D(K_r11[7]), .CK(n353), .Q(K_r12[7]) );
  DFFQX1 \K_r1_reg[6]  ( .D(K_r0[6]), .CK(n368), .Q(K_r1[6]) );
  DFFQX1 \K_r12_reg[6]  ( .D(K_r11[6]), .CK(n341), .Q(K_r12[6]) );
  DFFQX1 \K_r4_reg[5]  ( .D(K_r3[5]), .CK(n376), .Q(K_r4[5]) );
  DFFQX1 \K_r5_reg[5]  ( .D(K_r4[5]), .CK(n359), .Q(K_r5[5]) );
  DFFQX1 \K_r6_reg[5]  ( .D(K_r5[5]), .CK(n360), .Q(K_r6[5]) );
  DFFQX1 \K_r7_reg[5]  ( .D(K_r6[5]), .CK(n361), .Q(K_r7[5]) );
  DFFQX1 \K_r8_reg[5]  ( .D(K_r7[5]), .CK(n366), .Q(K_r8[5]) );
  DFFQX1 \K_r9_reg[5]  ( .D(K_r8[5]), .CK(n364), .Q(K_r9[5]) );
  DFFQX1 \K_r0_reg[4]  ( .D(K[4]), .CK(n347), .Q(K_r0[4]) );
  DFFQX1 \K_r2_reg[4]  ( .D(K_r1[4]), .CK(n348), .Q(K_r2[4]) );
  DFFQX1 \K_r3_reg[4]  ( .D(K_r2[4]), .CK(n349), .Q(K_r3[4]) );
  DFFQX1 \K_r10_reg[4]  ( .D(K_r9[4]), .CK(n354), .Q(K_r10[4]) );
  DFFQX1 \K_r11_reg[4]  ( .D(K_r10[4]), .CK(n355), .Q(K_r11[4]) );
  DFFQX1 \K_r13_reg[4]  ( .D(K_r12[4]), .CK(n356), .Q(K_r13[4]) );
  DFFQX1 \K_r0_reg[2]  ( .D(K[2]), .CK(n373), .Q(K_r0[2]) );
  DFFQX1 \K_r13_reg[2]  ( .D(K_r12[2]), .CK(n350), .Q(K_r13[2]) );
  DFFQX1 \K_r4_reg[0]  ( .D(K_r3[0]), .CK(n344), .Q(K_r4[0]) );
  DFFQX1 \K_r6_reg[0]  ( .D(K_r5[0]), .CK(n345), .Q(K_r6[0]) );
  DFFQX1 \K_r7_reg[0]  ( .D(K_r6[0]), .CK(n279), .Q(K_r7[0]) );
  DFFQX1 \K_r9_reg[0]  ( .D(K_r8[0]), .CK(n279), .Q(K_r9[0]) );
  DFFQX1 \K_r0_reg[55]  ( .D(K[55]), .CK(n341), .Q(K_r0[55]) );
  DFFQX1 \K_r1_reg[54]  ( .D(K_r0[54]), .CK(n339), .Q(K_r1[54]) );
  DFFQX1 \K_r12_reg[54]  ( .D(K_r11[54]), .CK(n338), .Q(K_r12[54]) );
  DFFQX1 \K_r1_reg[53]  ( .D(K_r0[53]), .CK(n338), .Q(K_r1[53]) );
  DFFQX1 \K_r12_reg[53]  ( .D(K_r11[53]), .CK(n336), .Q(K_r12[53]) );
  DFFQX1 \K_r1_reg[51]  ( .D(K_r0[51]), .CK(n334), .Q(K_r1[51]) );
  DFFQX1 \K_r12_reg[51]  ( .D(K_r11[51]), .CK(n333), .Q(K_r12[51]) );
  DFFQX1 \K_r1_reg[49]  ( .D(K_r0[49]), .CK(n331), .Q(K_r1[49]) );
  DFFQX1 \K_r12_reg[49]  ( .D(K_r11[49]), .CK(n330), .Q(K_r12[49]) );
  DFFQX1 \K_r1_reg[48]  ( .D(K_r0[48]), .CK(n330), .Q(K_r1[48]) );
  DFFQX1 \K_r12_reg[48]  ( .D(K_r11[48]), .CK(n329), .Q(K_r12[48]) );
  DFFQX1 \K_r1_reg[46]  ( .D(K_r0[46]), .CK(n327), .Q(K_r1[46]) );
  DFFQX1 \K_r12_reg[46]  ( .D(K_r11[46]), .CK(n325), .Q(K_r12[46]) );
  DFFQX1 \K_r1_reg[45]  ( .D(K_r0[45]), .CK(n325), .Q(K_r1[45]) );
  DFFQX1 \K_r12_reg[45]  ( .D(K_r11[45]), .CK(n324), .Q(K_r12[45]) );
  DFFQX1 \K_r1_reg[43]  ( .D(K_r0[43]), .CK(n322), .Q(K_r1[43]) );
  DFFQX1 \K_r12_reg[43]  ( .D(K_r11[43]), .CK(n321), .Q(K_r12[43]) );
  DFFQX1 \K_r1_reg[40]  ( .D(K_r0[40]), .CK(n317), .Q(K_r1[40]) );
  DFFQX1 \K_r12_reg[40]  ( .D(K_r11[40]), .CK(n316), .Q(K_r12[40]) );
  DFFQX1 \K_r1_reg[37]  ( .D(K_r0[37]), .CK(n313), .Q(K_r1[37]) );
  DFFQX1 \K_r12_reg[37]  ( .D(K_r11[37]), .CK(n311), .Q(K_r12[37]) );
  DFFQX1 \K_r1_reg[35]  ( .D(K_r0[35]), .CK(n310), .Q(K_r1[35]) );
  DFFQX1 \K_r12_reg[35]  ( .D(K_r11[35]), .CK(n308), .Q(K_r12[35]) );
  DFFQX1 \K_r1_reg[32]  ( .D(K_r0[32]), .CK(n305), .Q(K_r1[32]) );
  DFFQX1 \K_r12_reg[32]  ( .D(K_r11[32]), .CK(n304), .Q(K_r12[32]) );
  DFFQX1 \K_r1_reg[29]  ( .D(K_r0[29]), .CK(n300), .Q(K_r1[29]) );
  DFFQX1 \K_r12_reg[29]  ( .D(K_r11[29]), .CK(n299), .Q(K_r12[29]) );
  DFFQX1 \K_r1_reg[27]  ( .D(K_r0[27]), .CK(n297), .Q(K_r1[27]) );
  DFFQX1 \K_r12_reg[27]  ( .D(K_r11[27]), .CK(n296), .Q(K_r12[27]) );
  DFFQX1 \K_r1_reg[24]  ( .D(K_r0[24]), .CK(n292), .Q(K_r1[24]) );
  DFFQX1 \K_r12_reg[24]  ( .D(K_r11[24]), .CK(n291), .Q(K_r12[24]) );
  DFFQX1 \K_r1_reg[23]  ( .D(K_r0[23]), .CK(n291), .Q(K_r1[23]) );
  DFFQX1 \K_r12_reg[23]  ( .D(K_r11[23]), .CK(n290), .Q(K_r12[23]) );
  DFFQX1 \K_r1_reg[20]  ( .D(K_r0[20]), .CK(n286), .Q(K_r1[20]) );
  DFFQX1 \K_r12_reg[20]  ( .D(K_r11[20]), .CK(n285), .Q(K_r12[20]) );
  DFFQX1 \K_r1_reg[19]  ( .D(K_r0[19]), .CK(n285), .Q(K_r1[19]) );
  DFFQX1 \K_r12_reg[19]  ( .D(K_r11[19]), .CK(n283), .Q(K_r12[19]) );
  DFFQX1 \K_r1_reg[14]  ( .D(K_r0[14]), .CK(n370), .Q(K_r1[14]) );
  DFFQX1 \K_r12_reg[14]  ( .D(K_r11[14]), .CK(n366), .Q(K_r12[14]) );
  DFFQX1 \K_r1_reg[13]  ( .D(K_r0[13]), .CK(n368), .Q(K_r1[13]) );
  DFFQX1 \K_r12_reg[13]  ( .D(K_r11[13]), .CK(n348), .Q(K_r12[13]) );
  DFFQX1 \K_r1_reg[12]  ( .D(K_r0[12]), .CK(n349), .Q(K_r1[12]) );
  DFFQX1 \K_r12_reg[12]  ( .D(K_r11[12]), .CK(n363), .Q(K_r12[12]) );
  DFFQX1 \K_r1_reg[11]  ( .D(K_r0[11]), .CK(n368), .Q(K_r1[11]) );
  DFFQX1 \K_r12_reg[11]  ( .D(K_r11[11]), .CK(n349), .Q(K_r12[11]) );
  DFFQX1 \K_r1_reg[8]  ( .D(K_r0[8]), .CK(n352), .Q(K_r1[8]) );
  DFFQX1 \K_r12_reg[8]  ( .D(K_r11[8]), .CK(n359), .Q(K_r12[8]) );
  DFFQX1 \K_r1_reg[5]  ( .D(K_r0[5]), .CK(n342), .Q(K_r1[5]) );
  DFFQX1 \K_r12_reg[5]  ( .D(K_r11[5]), .CK(n360), .Q(K_r12[5]) );
  DFFQX1 \K_r1_reg[4]  ( .D(K_r0[4]), .CK(n370), .Q(K_r1[4]) );
  DFFQX1 \K_r12_reg[4]  ( .D(K_r11[4]), .CK(n357), .Q(K_r12[4]) );
  DFFQX1 \K_r1_reg[3]  ( .D(K_r0[3]), .CK(n358), .Q(K_r1[3]) );
  DFFQX1 \K_r12_reg[3]  ( .D(K_r11[3]), .CK(n373), .Q(K_r12[3]) );
  DFFQX1 \K_r1_reg[2]  ( .D(K_r0[2]), .CK(n371), .Q(K_r1[2]) );
  DFFQX1 \K_r12_reg[2]  ( .D(K_r11[2]), .CK(n351), .Q(K_r12[2]) );
  DFFQX1 \K_r1_reg[0]  ( .D(K_r0[0]), .CK(n346), .Q(K_r1[0]) );
  DFFQX1 \K_r12_reg[0]  ( .D(K_r11[0]), .CK(n279), .Q(K_r12[0]) );
  DFFQX1 \K_r14_reg[52]  ( .D(K_r13[52]), .CK(n278), .Q(K_r14[52]) );
  DFFQX1 \K_r14_reg[25]  ( .D(K_r13[25]), .CK(n275), .Q(K_r14[25]) );
  DFFQX1 \K_r14_reg[22]  ( .D(K_r13[22]), .CK(n275), .Q(K_r14[22]) );
  DFFQX1 \K_r14_reg[19]  ( .D(K_r13[19]), .CK(n275), .Q(K_r14[19]) );
  DFFQX1 \K_r14_reg[17]  ( .D(K_r13[17]), .CK(n274), .Q(K_r14[17]) );
  DFFQX1 \K_r14_reg[55]  ( .D(K_r13[55]), .CK(n279), .Q(K_r14[55]) );
  DFFQX1 \K_r14_reg[54]  ( .D(K_r13[54]), .CK(n279), .Q(K_r14[54]) );
  DFFQX1 \K_r14_reg[51]  ( .D(K_r13[51]), .CK(n278), .Q(K_r14[51]) );
  DFFQX1 \K_r14_reg[48]  ( .D(K_r13[48]), .CK(n278), .Q(K_r14[48]) );
  DFFQX1 \K_r14_reg[47]  ( .D(K_r13[47]), .CK(n278), .Q(K_r14[47]) );
  DFFQX1 \K_r14_reg[44]  ( .D(K_r13[44]), .CK(n277), .Q(K_r14[44]) );
  DFFQX1 \K_r14_reg[41]  ( .D(K_r13[41]), .CK(n277), .Q(K_r14[41]) );
  DFFQX1 \K_r14_reg[37]  ( .D(K_r13[37]), .CK(n277), .Q(K_r14[37]) );
  DFFQX1 \K_r14_reg[36]  ( .D(K_r13[36]), .CK(n277), .Q(K_r14[36]) );
  DFFQX1 \K_r14_reg[35]  ( .D(K_r13[35]), .CK(n276), .Q(K_r14[35]) );
  DFFQX1 \K_r14_reg[34]  ( .D(K_r13[34]), .CK(n276), .Q(K_r14[34]) );
  DFFQX1 \K_r14_reg[33]  ( .D(K_r13[33]), .CK(n276), .Q(K_r14[33]) );
  DFFQX1 \K_r14_reg[31]  ( .D(K_r13[31]), .CK(n276), .Q(K_r14[31]) );
  DFFQX1 \K_r14_reg[28]  ( .D(K_r13[28]), .CK(n276), .Q(K_r14[28]) );
  DFFQX1 \K_r14_reg[26]  ( .D(K_r13[26]), .CK(n275), .Q(K_r14[26]) );
  DFFQX1 \K_r14_reg[24]  ( .D(K_r13[24]), .CK(n275), .Q(K_r14[24]) );
  DFFQX1 \K_r14_reg[23]  ( .D(K_r13[23]), .CK(n275), .Q(K_r14[23]) );
  DFFQX1 \K_r14_reg[21]  ( .D(K_r13[21]), .CK(n275), .Q(K_r14[21]) );
  DFFQX1 \K_r14_reg[20]  ( .D(K_r13[20]), .CK(n275), .Q(K_r14[20]) );
  DFFQX1 \K_r14_reg[16]  ( .D(K_r13[16]), .CK(n274), .Q(K_r14[16]) );
  DFFQX1 \K_r14_reg[13]  ( .D(K_r13[13]), .CK(n274), .Q(K_r14[13]) );
  DFFQX1 \K_r14_reg[9]  ( .D(K_r13[9]), .CK(n274), .Q(K_r14[9]) );
  DFFQX1 \K_r14_reg[7]  ( .D(K_r13[7]), .CK(n273), .Q(K_r14[7]) );
  DFFQX1 \K_r14_reg[6]  ( .D(K_r13[6]), .CK(n273), .Q(K_r14[6]) );
  DFFQX1 \K_r14_reg[4]  ( .D(K_r13[4]), .CK(n273), .Q(K_r14[4]) );
  DFFQX1 \K_r14_reg[2]  ( .D(K_r13[2]), .CK(n273), .Q(K_r14[2]) );
  DFFQX1 \K_r14_reg[0]  ( .D(K_r13[0]), .CK(n273), .Q(K_r14[0]) );
  DFFQX1 \K_r14_reg[53]  ( .D(K_r13[53]), .CK(n278), .Q(K_r14[53]) );
  DFFQX1 \K_r14_reg[40]  ( .D(K_r13[40]), .CK(n277), .Q(K_r14[40]) );
  DFFQX1 \K_r14_reg[32]  ( .D(K_r13[32]), .CK(n276), .Q(K_r14[32]) );
  DFFQX1 \K_r14_reg[30]  ( .D(K_r13[30]), .CK(n276), .Q(K_r14[30]) );
  DFFQX1 \K_r14_reg[29]  ( .D(K_r13[29]), .CK(n276), .Q(K_r14[29]) );
  DFFQX1 \K_r14_reg[27]  ( .D(K_r13[27]), .CK(n276), .Q(K_r14[27]) );
  DFFQX1 \K_r14_reg[14]  ( .D(K_r13[14]), .CK(n274), .Q(K_r14[14]) );
  DFFQX1 \K_r14_reg[1]  ( .D(K_r13[1]), .CK(n273), .Q(K_r14[1]) );
  DFFQX1 \K_r3_reg[53]  ( .D(K_r2[53]), .CK(n337), .Q(K_r3[53]) );
  DFFQX1 \K_r11_reg[51]  ( .D(K_r10[51]), .CK(n333), .Q(K_r11[51]) );
  DFFQX1 \K_r3_reg[50]  ( .D(K_r2[50]), .CK(n333), .Q(K_r3[50]) );
  DFFQX1 \K_r9_reg[50]  ( .D(K_r8[50]), .CK(n332), .Q(K_r9[50]) );
  DFFQX1 \K_r9_reg[46]  ( .D(K_r8[46]), .CK(n326), .Q(K_r9[46]) );
  DFFQX1 \K_r13_reg[46]  ( .D(K_r12[46]), .CK(n325), .Q(K_r13[46]) );
  DFFQX1 \K_r4_reg[43]  ( .D(K_r3[43]), .CK(n322), .Q(K_r4[43]) );
  DFFQX1 \K_r11_reg[43]  ( .D(K_r10[43]), .CK(n321), .Q(K_r11[43]) );
  DFFQX1 \K_r13_reg[43]  ( .D(K_r12[43]), .CK(n321), .Q(K_r13[43]) );
  DFFQX1 \K_r4_reg[42]  ( .D(K_r3[42]), .CK(n320), .Q(K_r4[42]) );
  DFFQX1 \K_r6_reg[41]  ( .D(K_r5[41]), .CK(n318), .Q(K_r6[41]) );
  DFFQX1 \K_r11_reg[40]  ( .D(K_r10[40]), .CK(n316), .Q(K_r11[40]) );
  DFFQX1 \K_r4_reg[39]  ( .D(K_r3[39]), .CK(n315), .Q(K_r4[39]) );
  DFFQX1 \K_r6_reg[38]  ( .D(K_r5[38]), .CK(n314), .Q(K_r6[38]) );
  DFFQX1 \K_r12_reg[38]  ( .D(K_r11[38]), .CK(n313), .Q(K_r12[38]) );
  DFFQX1 \K_r0_reg[37]  ( .D(K[37]), .CK(n313), .Q(K_r0[37]) );
  DFFQX1 \K_r2_reg[37]  ( .D(K_r1[37]), .CK(n313), .Q(K_r2[37]) );
  DFFQX1 \K_r6_reg[36]  ( .D(K_r5[36]), .CK(n311), .Q(K_r6[36]) );
  DFFQX1 \K_r8_reg[36]  ( .D(K_r7[36]), .CK(n310), .Q(K_r8[36]) );
  DFFQX1 \K_r6_reg[33]  ( .D(K_r5[33]), .CK(n306), .Q(K_r6[33]) );
  DFFQX1 \K_r2_reg[32]  ( .D(K_r1[32]), .CK(n305), .Q(K_r2[32]) );
  DFFQX1 \K_r1_reg[28]  ( .D(K_r0[28]), .CK(n299), .Q(K_r1[28]) );
  DFFQX1 \K_r3_reg[21]  ( .D(K_r2[21]), .CK(n288), .Q(K_r3[21]) );
  DFFQX1 \K_r3_reg[20]  ( .D(K_r2[20]), .CK(n286), .Q(K_r3[20]) );
  DFFQX1 \K_r5_reg[20]  ( .D(K_r4[20]), .CK(n286), .Q(K_r5[20]) );
  DFFQX1 \K_r7_reg[13]  ( .D(K_r6[13]), .CK(n356), .Q(K_r7[13]) );
  DFFQX1 \K_r4_reg[8]  ( .D(K_r3[8]), .CK(n347), .Q(K_r4[8]) );
  DFFQX1 \K_r10_reg[8]  ( .D(K_r9[8]), .CK(n348), .Q(K_r10[8]) );
  DFFQX1 \K_r10_reg[7]  ( .D(K_r9[7]), .CK(n364), .Q(K_r10[7]) );
  DFFQX1 \K_r7_reg[6]  ( .D(K_r6[6]), .CK(n356), .Q(K_r7[6]) );
  DFFQX1 \K_r2_reg[5]  ( .D(K_r1[5]), .CK(n343), .Q(K_r2[5]) );
  DFFQX1 \K_r8_reg[3]  ( .D(K_r7[3]), .CK(n374), .Q(K_r8[3]) );
  DFFQX1 \K_r3_reg[55]  ( .D(K_r2[55]), .CK(n340), .Q(K_r3[55]) );
  DFFQX1 \K_r5_reg[55]  ( .D(K_r4[55]), .CK(n340), .Q(K_r5[55]) );
  DFFQX1 \K_r8_reg[55]  ( .D(K_r7[55]), .CK(n340), .Q(K_r8[55]) );
  DFFQX1 \K_r10_reg[55]  ( .D(K_r9[55]), .CK(n340), .Q(K_r10[55]) );
  DFFQX1 \K_r0_reg[54]  ( .D(K[54]), .CK(n339), .Q(K_r0[54]) );
  DFFQX1 \K_r3_reg[54]  ( .D(K_r2[54]), .CK(n339), .Q(K_r3[54]) );
  DFFQX1 \K_r6_reg[54]  ( .D(K_r5[54]), .CK(n339), .Q(K_r6[54]) );
  DFFQX1 \K_r7_reg[54]  ( .D(K_r6[54]), .CK(n338), .Q(K_r7[54]) );
  DFFQX1 \K_r10_reg[54]  ( .D(K_r9[54]), .CK(n338), .Q(K_r10[54]) );
  DFFQX1 \K_r13_reg[54]  ( .D(K_r12[54]), .CK(n338), .Q(K_r13[54]) );
  DFFQX1 \K_r8_reg[53]  ( .D(K_r7[53]), .CK(n337), .Q(K_r8[53]) );
  DFFQX1 \K_r10_reg[53]  ( .D(K_r9[53]), .CK(n337), .Q(K_r10[53]) );
  DFFQX1 \K_r2_reg[52]  ( .D(K_r1[52]), .CK(n336), .Q(K_r2[52]) );
  DFFQX1 \K_r4_reg[52]  ( .D(K_r3[52]), .CK(n336), .Q(K_r4[52]) );
  DFFQX1 \K_r5_reg[52]  ( .D(K_r4[52]), .CK(n336), .Q(K_r5[52]) );
  DFFQX1 \K_r6_reg[52]  ( .D(K_r5[52]), .CK(n335), .Q(K_r6[52]) );
  DFFQX1 \K_r8_reg[52]  ( .D(K_r7[52]), .CK(n335), .Q(K_r8[52]) );
  DFFQX1 \K_r11_reg[52]  ( .D(K_r10[52]), .CK(n335), .Q(K_r11[52]) );
  DFFQX1 \K_r0_reg[51]  ( .D(K[51]), .CK(n335), .Q(K_r0[51]) );
  DFFQX1 \K_r2_reg[51]  ( .D(K_r1[51]), .CK(n334), .Q(K_r2[51]) );
  DFFQX1 \K_r3_reg[51]  ( .D(K_r2[51]), .CK(n334), .Q(K_r3[51]) );
  DFFQX1 \K_r4_reg[51]  ( .D(K_r3[51]), .CK(n334), .Q(K_r4[51]) );
  DFFQX1 \K_r9_reg[51]  ( .D(K_r8[51]), .CK(n334), .Q(K_r9[51]) );
  DFFQX1 \K_r10_reg[51]  ( .D(K_r9[51]), .CK(n333), .Q(K_r10[51]) );
  DFFQX1 \K_r13_reg[51]  ( .D(K_r12[51]), .CK(n333), .Q(K_r13[51]) );
  DFFQX1 \K_r0_reg[50]  ( .D(K[50]), .CK(n333), .Q(K_r0[50]) );
  DFFQX1 \K_r5_reg[50]  ( .D(K_r4[50]), .CK(n332), .Q(K_r5[50]) );
  DFFQX1 \K_r6_reg[50]  ( .D(K_r5[50]), .CK(n332), .Q(K_r6[50]) );
  DFFQX1 \K_r7_reg[50]  ( .D(K_r6[50]), .CK(n332), .Q(K_r7[50]) );
  DFFQX1 \K_r8_reg[50]  ( .D(K_r7[50]), .CK(n332), .Q(K_r8[50]) );
  DFFQX1 \K_r10_reg[50]  ( .D(K_r9[50]), .CK(n332), .Q(K_r10[50]) );
  DFFQX1 \K_r13_reg[50]  ( .D(K_r12[50]), .CK(n332), .Q(K_r13[50]) );
  DFFQX1 \K_r0_reg[49]  ( .D(K[49]), .CK(n331), .Q(K_r0[49]) );
  DFFQX1 \K_r2_reg[49]  ( .D(K_r1[49]), .CK(n331), .Q(K_r2[49]) );
  DFFQX1 \K_r5_reg[49]  ( .D(K_r4[49]), .CK(n331), .Q(K_r5[49]) );
  DFFQX1 \K_r6_reg[49]  ( .D(K_r5[49]), .CK(n331), .Q(K_r6[49]) );
  DFFQX1 \K_r7_reg[49]  ( .D(K_r6[49]), .CK(n331), .Q(K_r7[49]) );
  DFFQX1 \K_r8_reg[49]  ( .D(K_r7[49]), .CK(n331), .Q(K_r8[49]) );
  DFFQX1 \K_r11_reg[49]  ( .D(K_r10[49]), .CK(n330), .Q(K_r11[49]) );
  DFFQX1 \K_r13_reg[49]  ( .D(K_r12[49]), .CK(n330), .Q(K_r13[49]) );
  DFFQX1 \K_r0_reg[48]  ( .D(K[48]), .CK(n330), .Q(K_r0[48]) );
  DFFQX1 \K_r2_reg[48]  ( .D(K_r1[48]), .CK(n330), .Q(K_r2[48]) );
  DFFQX1 \K_r3_reg[48]  ( .D(K_r2[48]), .CK(n330), .Q(K_r3[48]) );
  DFFQX1 \K_r10_reg[48]  ( .D(K_r9[48]), .CK(n329), .Q(K_r10[48]) );
  DFFQX1 \K_r11_reg[48]  ( .D(K_r10[48]), .CK(n329), .Q(K_r11[48]) );
  DFFQX1 \K_r13_reg[48]  ( .D(K_r12[48]), .CK(n328), .Q(K_r13[48]) );
  DFFQX1 \K_r0_reg[47]  ( .D(K[47]), .CK(n328), .Q(K_r0[47]) );
  DFFQX1 \K_r4_reg[47]  ( .D(K_r3[47]), .CK(n328), .Q(K_r4[47]) );
  DFFQX1 \K_r5_reg[47]  ( .D(K_r4[47]), .CK(n328), .Q(K_r5[47]) );
  DFFQX1 \K_r6_reg[47]  ( .D(K_r5[47]), .CK(n328), .Q(K_r6[47]) );
  DFFQX1 \K_r7_reg[47]  ( .D(K_r6[47]), .CK(n328), .Q(K_r7[47]) );
  DFFQX1 \K_r8_reg[47]  ( .D(K_r7[47]), .CK(n327), .Q(K_r8[47]) );
  DFFQX1 \K_r9_reg[47]  ( .D(K_r8[47]), .CK(n327), .Q(K_r9[47]) );
  DFFQX1 \K_r13_reg[47]  ( .D(K_r12[47]), .CK(n327), .Q(K_r13[47]) );
  DFFQX1 \K_r0_reg[46]  ( .D(K[46]), .CK(n327), .Q(K_r0[46]) );
  DFFQX1 \K_r2_reg[46]  ( .D(K_r1[46]), .CK(n327), .Q(K_r2[46]) );
  DFFQX1 \K_r3_reg[46]  ( .D(K_r2[46]), .CK(n326), .Q(K_r3[46]) );
  DFFQX1 \K_r4_reg[46]  ( .D(K_r3[46]), .CK(n326), .Q(K_r4[46]) );
  DFFQX1 \K_r8_reg[46]  ( .D(K_r7[46]), .CK(n326), .Q(K_r8[46]) );
  DFFQX1 \K_r10_reg[46]  ( .D(K_r9[46]), .CK(n326), .Q(K_r10[46]) );
  DFFQX1 \K_r11_reg[46]  ( .D(K_r10[46]), .CK(n326), .Q(K_r11[46]) );
  DFFQX1 \K_r4_reg[45]  ( .D(K_r3[45]), .CK(n325), .Q(K_r4[45]) );
  DFFQX1 \K_r7_reg[45]  ( .D(K_r6[45]), .CK(n324), .Q(K_r7[45]) );
  DFFQX1 \K_r9_reg[45]  ( .D(K_r8[45]), .CK(n324), .Q(K_r9[45]) );
  DFFQX1 \K_r13_reg[45]  ( .D(K_r12[45]), .CK(n324), .Q(K_r13[45]) );
  DFFQX1 \K_r0_reg[44]  ( .D(K[44]), .CK(n324), .Q(K_r0[44]) );
  DFFQX1 \K_r4_reg[44]  ( .D(K_r3[44]), .CK(n323), .Q(K_r4[44]) );
  DFFQX1 \K_r5_reg[44]  ( .D(K_r4[44]), .CK(n323), .Q(K_r5[44]) );
  DFFQX1 \K_r8_reg[44]  ( .D(K_r7[44]), .CK(n323), .Q(K_r8[44]) );
  DFFQX1 \K_r9_reg[44]  ( .D(K_r8[44]), .CK(n323), .Q(K_r9[44]) );
  DFFQX1 \K_r13_reg[44]  ( .D(K_r12[44]), .CK(n322), .Q(K_r13[44]) );
  DFFQX1 \K_r0_reg[43]  ( .D(K[43]), .CK(n322), .Q(K_r0[43]) );
  DFFQX1 \K_r2_reg[43]  ( .D(K_r1[43]), .CK(n322), .Q(K_r2[43]) );
  DFFQX1 \K_r6_reg[43]  ( .D(K_r5[43]), .CK(n321), .Q(K_r6[43]) );
  DFFQX1 \K_r7_reg[43]  ( .D(K_r6[43]), .CK(n321), .Q(K_r7[43]) );
  DFFQX1 \K_r9_reg[43]  ( .D(K_r8[43]), .CK(n321), .Q(K_r9[43]) );
  DFFQX1 \K_r2_reg[42]  ( .D(K_r1[42]), .CK(n320), .Q(K_r2[42]) );
  DFFQX1 \K_r3_reg[42]  ( .D(K_r2[42]), .CK(n320), .Q(K_r3[42]) );
  DFFQX1 \K_r5_reg[42]  ( .D(K_r4[42]), .CK(n320), .Q(K_r5[42]) );
  DFFQX1 \K_r8_reg[42]  ( .D(K_r7[42]), .CK(n320), .Q(K_r8[42]) );
  DFFQX1 \K_r10_reg[42]  ( .D(K_r9[42]), .CK(n319), .Q(K_r10[42]) );
  DFFQX1 \K_r11_reg[42]  ( .D(K_r10[42]), .CK(n319), .Q(K_r11[42]) );
  DFFQX1 \K_r0_reg[41]  ( .D(K[41]), .CK(n319), .Q(K_r0[41]) );
  DFFQX1 \K_r2_reg[41]  ( .D(K_r1[41]), .CK(n319), .Q(K_r2[41]) );
  DFFQX1 \K_r3_reg[41]  ( .D(K_r2[41]), .CK(n319), .Q(K_r3[41]) );
  DFFQX1 \K_r4_reg[41]  ( .D(K_r3[41]), .CK(n319), .Q(K_r4[41]) );
  DFFQX1 \K_r7_reg[41]  ( .D(K_r6[41]), .CK(n318), .Q(K_r7[41]) );
  DFFQX1 \K_r9_reg[41]  ( .D(K_r8[41]), .CK(n318), .Q(K_r9[41]) );
  DFFQX1 \K_r10_reg[41]  ( .D(K_r9[41]), .CK(n318), .Q(K_r10[41]) );
  DFFQX1 \K_r11_reg[41]  ( .D(K_r10[41]), .CK(n318), .Q(K_r11[41]) );
  DFFQX1 \K_r13_reg[41]  ( .D(K_r12[41]), .CK(n318), .Q(K_r13[41]) );
  DFFQX1 \K_r2_reg[40]  ( .D(K_r1[40]), .CK(n317), .Q(K_r2[40]) );
  DFFQX1 \K_r3_reg[40]  ( .D(K_r2[40]), .CK(n317), .Q(K_r3[40]) );
  DFFQX1 \K_r4_reg[40]  ( .D(K_r3[40]), .CK(n317), .Q(K_r4[40]) );
  DFFQX1 \K_r6_reg[40]  ( .D(K_r5[40]), .CK(n317), .Q(K_r6[40]) );
  DFFQX1 \K_r7_reg[40]  ( .D(K_r6[40]), .CK(n317), .Q(K_r7[40]) );
  DFFQX1 \K_r9_reg[40]  ( .D(K_r8[40]), .CK(n316), .Q(K_r9[40]) );
  DFFQX1 \K_r10_reg[40]  ( .D(K_r9[40]), .CK(n316), .Q(K_r10[40]) );
  DFFQX1 \K_r2_reg[39]  ( .D(K_r1[39]), .CK(n316), .Q(K_r2[39]) );
  DFFQX1 \K_r6_reg[39]  ( .D(K_r5[39]), .CK(n315), .Q(K_r6[39]) );
  DFFQX1 \K_r7_reg[39]  ( .D(K_r6[39]), .CK(n315), .Q(K_r7[39]) );
  DFFQX1 \K_r9_reg[39]  ( .D(K_r8[39]), .CK(n315), .Q(K_r9[39]) );
  DFFQX1 \K_r11_reg[39]  ( .D(K_r10[39]), .CK(n315), .Q(K_r11[39]) );
  DFFQX1 \K_r0_reg[38]  ( .D(K[38]), .CK(n314), .Q(K_r0[38]) );
  DFFQX1 \K_r2_reg[38]  ( .D(K_r1[38]), .CK(n314), .Q(K_r2[38]) );
  DFFQX1 \K_r3_reg[38]  ( .D(K_r2[38]), .CK(n314), .Q(K_r3[38]) );
  DFFQX1 \K_r5_reg[38]  ( .D(K_r4[38]), .CK(n314), .Q(K_r5[38]) );
  DFFQX1 \K_r7_reg[38]  ( .D(K_r6[38]), .CK(n314), .Q(K_r7[38]) );
  DFFQX1 \K_r8_reg[38]  ( .D(K_r7[38]), .CK(n313), .Q(K_r8[38]) );
  DFFQX1 \K_r10_reg[38]  ( .D(K_r9[38]), .CK(n313), .Q(K_r10[38]) );
  DFFQX1 \K_r11_reg[38]  ( .D(K_r10[38]), .CK(n313), .Q(K_r11[38]) );
  DFFQX1 \K_r13_reg[38]  ( .D(K_r12[38]), .CK(n313), .Q(K_r13[38]) );
  DFFQX1 \K_r3_reg[37]  ( .D(K_r2[37]), .CK(n312), .Q(K_r3[37]) );
  DFFQX1 \K_r4_reg[37]  ( .D(K_r3[37]), .CK(n312), .Q(K_r4[37]) );
  DFFQX1 \K_r9_reg[37]  ( .D(K_r8[37]), .CK(n312), .Q(K_r9[37]) );
  DFFQX1 \K_r10_reg[37]  ( .D(K_r9[37]), .CK(n312), .Q(K_r10[37]) );
  DFFQX1 \K_r11_reg[37]  ( .D(K_r10[37]), .CK(n312), .Q(K_r11[37]) );
  DFFQX1 \K_r13_reg[37]  ( .D(K_r12[37]), .CK(n311), .Q(K_r13[37]) );
  DFFQX1 \K_r2_reg[36]  ( .D(K_r1[36]), .CK(n311), .Q(K_r2[36]) );
  DFFQX1 \K_r3_reg[36]  ( .D(K_r2[36]), .CK(n311), .Q(K_r3[36]) );
  DFFQX1 \K_r4_reg[36]  ( .D(K_r3[36]), .CK(n311), .Q(K_r4[36]) );
  DFFQX1 \K_r7_reg[36]  ( .D(K_r6[36]), .CK(n310), .Q(K_r7[36]) );
  DFFQX1 \K_r9_reg[36]  ( .D(K_r8[36]), .CK(n310), .Q(K_r9[36]) );
  DFFQX1 \K_r10_reg[36]  ( .D(K_r9[36]), .CK(n310), .Q(K_r10[36]) );
  DFFQX1 \K_r11_reg[36]  ( .D(K_r10[36]), .CK(n310), .Q(K_r11[36]) );
  DFFQX1 \K_r2_reg[35]  ( .D(K_r1[35]), .CK(n309), .Q(K_r2[35]) );
  DFFQX1 \K_r5_reg[35]  ( .D(K_r4[35]), .CK(n309), .Q(K_r5[35]) );
  DFFQX1 \K_r6_reg[35]  ( .D(K_r5[35]), .CK(n309), .Q(K_r6[35]) );
  DFFQX1 \K_r7_reg[35]  ( .D(K_r6[35]), .CK(n309), .Q(K_r7[35]) );
  DFFQX1 \K_r8_reg[35]  ( .D(K_r7[35]), .CK(n309), .Q(K_r8[35]) );
  DFFQX1 \K_r11_reg[35]  ( .D(K_r10[35]), .CK(n308), .Q(K_r11[35]) );
  DFFQX1 \K_r1_reg[34]  ( .D(K_r0[34]), .CK(n308), .Q(K_r1[34]) );
  DFFQX1 \K_r2_reg[34]  ( .D(K_r1[34]), .CK(n308), .Q(K_r2[34]) );
  DFFQX1 \K_r4_reg[34]  ( .D(K_r3[34]), .CK(n308), .Q(K_r4[34]) );
  DFFQX1 \K_r5_reg[34]  ( .D(K_r4[34]), .CK(n308), .Q(K_r5[34]) );
  DFFQX1 \K_r8_reg[34]  ( .D(K_r7[34]), .CK(n307), .Q(K_r8[34]) );
  DFFQX1 \K_r9_reg[34]  ( .D(K_r8[34]), .CK(n307), .Q(K_r9[34]) );
  DFFQX1 \K_r11_reg[34]  ( .D(K_r10[34]), .CK(n307), .Q(K_r11[34]) );
  DFFQX1 \K_r0_reg[33]  ( .D(K[33]), .CK(n307), .Q(K_r0[33]) );
  DFFQX1 \K_r3_reg[33]  ( .D(K_r2[33]), .CK(n306), .Q(K_r3[33]) );
  DFFQX1 \K_r5_reg[33]  ( .D(K_r4[33]), .CK(n306), .Q(K_r5[33]) );
  DFFQX1 \K_r7_reg[33]  ( .D(K_r6[33]), .CK(n306), .Q(K_r7[33]) );
  DFFQX1 \K_r8_reg[33]  ( .D(K_r7[33]), .CK(n306), .Q(K_r8[33]) );
  DFFQX1 \K_r13_reg[33]  ( .D(K_r12[33]), .CK(n305), .Q(K_r13[33]) );
  DFFQX1 \K_r3_reg[32]  ( .D(K_r2[32]), .CK(n305), .Q(K_r3[32]) );
  DFFQX1 \K_r6_reg[32]  ( .D(K_r5[32]), .CK(n304), .Q(K_r6[32]) );
  DFFQX1 \K_r7_reg[32]  ( .D(K_r6[32]), .CK(n304), .Q(K_r7[32]) );
  DFFQX1 \K_r9_reg[32]  ( .D(K_r8[32]), .CK(n304), .Q(K_r9[32]) );
  DFFQX1 \K_r10_reg[32]  ( .D(K_r9[32]), .CK(n304), .Q(K_r10[32]) );
  DFFQX1 \K_r11_reg[32]  ( .D(K_r10[32]), .CK(n304), .Q(K_r11[32]) );
  DFFQX1 \K_r2_reg[31]  ( .D(K_r1[31]), .CK(n303), .Q(K_r2[31]) );
  DFFQX1 \K_r3_reg[31]  ( .D(K_r2[31]), .CK(n303), .Q(K_r3[31]) );
  DFFQX1 \K_r5_reg[31]  ( .D(K_r4[31]), .CK(n303), .Q(K_r5[31]) );
  DFFQX1 \K_r8_reg[31]  ( .D(K_r7[31]), .CK(n303), .Q(K_r8[31]) );
  DFFQX1 \K_r10_reg[31]  ( .D(K_r9[31]), .CK(n302), .Q(K_r10[31]) );
  DFFQX1 \K_r11_reg[31]  ( .D(K_r10[31]), .CK(n302), .Q(K_r11[31]) );
  DFFQX1 \K_r12_reg[31]  ( .D(K_r11[31]), .CK(n302), .Q(K_r12[31]) );
  DFFQX1 \K_r0_reg[30]  ( .D(K[30]), .CK(n302), .Q(K_r0[30]) );
  DFFQX1 \K_r1_reg[30]  ( .D(K_r0[30]), .CK(n302), .Q(K_r1[30]) );
  DFFQX1 \K_r4_reg[30]  ( .D(K_r3[30]), .CK(n301), .Q(K_r4[30]) );
  DFFQX1 \K_r5_reg[30]  ( .D(K_r4[30]), .CK(n301), .Q(K_r5[30]) );
  DFFQX1 \K_r8_reg[30]  ( .D(K_r7[30]), .CK(n301), .Q(K_r8[30]) );
  DFFQX1 \K_r9_reg[30]  ( .D(K_r8[30]), .CK(n301), .Q(K_r9[30]) );
  DFFQX1 \K_r12_reg[30]  ( .D(K_r11[30]), .CK(n301), .Q(K_r12[30]) );
  DFFQX1 \K_r13_reg[30]  ( .D(K_r12[30]), .CK(n300), .Q(K_r13[30]) );
  DFFQX1 \K_r0_reg[29]  ( .D(K[29]), .CK(n300), .Q(K_r0[29]) );
  DFFQX1 \K_r3_reg[29]  ( .D(K_r2[29]), .CK(n300), .Q(K_r3[29]) );
  DFFQX1 \K_r5_reg[29]  ( .D(K_r4[29]), .CK(n300), .Q(K_r5[29]) );
  DFFQX1 \K_r8_reg[29]  ( .D(K_r7[29]), .CK(n299), .Q(K_r8[29]) );
  DFFQX1 \K_r10_reg[29]  ( .D(K_r9[29]), .CK(n299), .Q(K_r10[29]) );
  DFFQX1 \K_r13_reg[29]  ( .D(K_r12[29]), .CK(n299), .Q(K_r13[29]) );
  DFFQX1 \K_r0_reg[28]  ( .D(K[28]), .CK(n299), .Q(K_r0[28]) );
  DFFQX1 \K_r3_reg[28]  ( .D(K_r2[28]), .CK(n298), .Q(K_r3[28]) );
  DFFQX1 \K_r4_reg[28]  ( .D(K_r3[28]), .CK(n298), .Q(K_r4[28]) );
  DFFQX1 \K_r5_reg[28]  ( .D(K_r4[28]), .CK(n298), .Q(K_r5[28]) );
  DFFQX1 \K_r6_reg[28]  ( .D(K_r5[28]), .CK(n298), .Q(K_r6[28]) );
  DFFQX1 \K_r7_reg[28]  ( .D(K_r6[28]), .CK(n298), .Q(K_r7[28]) );
  DFFQX1 \K_r8_reg[28]  ( .D(K_r7[28]), .CK(n298), .Q(K_r8[28]) );
  DFFQX1 \K_r9_reg[28]  ( .D(K_r8[28]), .CK(n298), .Q(K_r9[28]) );
  DFFQX1 \K_r10_reg[28]  ( .D(K_r9[28]), .CK(n298), .Q(K_r10[28]) );
  DFFQX1 \K_r13_reg[28]  ( .D(K_r12[28]), .CK(n297), .Q(K_r13[28]) );
  DFFQX1 \K_r0_reg[27]  ( .D(K[27]), .CK(n297), .Q(K_r0[27]) );
  DFFQX1 \K_r3_reg[27]  ( .D(K_r2[27]), .CK(n297), .Q(K_r3[27]) );
  DFFQX1 \K_r5_reg[27]  ( .D(K_r4[27]), .CK(n297), .Q(K_r5[27]) );
  DFFQX1 \K_r8_reg[27]  ( .D(K_r7[27]), .CK(n296), .Q(K_r8[27]) );
  DFFQX1 \K_r10_reg[27]  ( .D(K_r9[27]), .CK(n296), .Q(K_r10[27]) );
  DFFQX1 \K_r13_reg[27]  ( .D(K_r12[27]), .CK(n296), .Q(K_r13[27]) );
  DFFQX1 \K_r0_reg[26]  ( .D(K[26]), .CK(n296), .Q(K_r0[26]) );
  DFFQX1 \K_r3_reg[26]  ( .D(K_r2[26]), .CK(n295), .Q(K_r3[26]) );
  DFFQX1 \K_r4_reg[26]  ( .D(K_r3[26]), .CK(n295), .Q(K_r4[26]) );
  DFFQX1 \K_r5_reg[26]  ( .D(K_r4[26]), .CK(n295), .Q(K_r5[26]) );
  DFFQX1 \K_r8_reg[26]  ( .D(K_r7[26]), .CK(n295), .Q(K_r8[26]) );
  DFFQX1 \K_r9_reg[26]  ( .D(K_r8[26]), .CK(n295), .Q(K_r9[26]) );
  DFFQX1 \K_r10_reg[26]  ( .D(K_r9[26]), .CK(n295), .Q(K_r10[26]) );
  DFFQX1 \K_r12_reg[26]  ( .D(K_r11[26]), .CK(n294), .Q(K_r12[26]) );
  DFFQX1 \K_r13_reg[26]  ( .D(K_r12[26]), .CK(n294), .Q(K_r13[26]) );
  DFFQX1 \K_r3_reg[25]  ( .D(K_r2[25]), .CK(n294), .Q(K_r3[25]) );
  DFFQX1 \K_r4_reg[25]  ( .D(K_r3[25]), .CK(n294), .Q(K_r4[25]) );
  DFFQX1 \K_r5_reg[25]  ( .D(K_r4[25]), .CK(n294), .Q(K_r5[25]) );
  DFFQX1 \K_r6_reg[25]  ( .D(K_r5[25]), .CK(n293), .Q(K_r6[25]) );
  DFFQX1 \K_r7_reg[25]  ( .D(K_r6[25]), .CK(n293), .Q(K_r7[25]) );
  DFFQX1 \K_r8_reg[25]  ( .D(K_r7[25]), .CK(n293), .Q(K_r8[25]) );
  DFFQX1 \K_r9_reg[25]  ( .D(K_r8[25]), .CK(n293), .Q(K_r9[25]) );
  DFFQX1 \K_r10_reg[25]  ( .D(K_r9[25]), .CK(n293), .Q(K_r10[25]) );
  DFFQX1 \K_r0_reg[24]  ( .D(K[24]), .CK(n293), .Q(K_r0[24]) );
  DFFQX1 \K_r5_reg[24]  ( .D(K_r4[24]), .CK(n292), .Q(K_r5[24]) );
  DFFQX1 \K_r10_reg[24]  ( .D(K_r9[24]), .CK(n291), .Q(K_r10[24]) );
  DFFQX1 \K_r13_reg[24]  ( .D(K_r12[24]), .CK(n291), .Q(K_r13[24]) );
  DFFQX1 \K_r0_reg[23]  ( .D(K[23]), .CK(n291), .Q(K_r0[23]) );
  DFFQX1 \K_r2_reg[23]  ( .D(K_r1[23]), .CK(n291), .Q(K_r2[23]) );
  DFFQX1 \K_r3_reg[23]  ( .D(K_r2[23]), .CK(n291), .Q(K_r3[23]) );
  DFFQX1 \K_r5_reg[23]  ( .D(K_r4[23]), .CK(n290), .Q(K_r5[23]) );
  DFFQX1 \K_r6_reg[23]  ( .D(K_r5[23]), .CK(n290), .Q(K_r6[23]) );
  DFFQX1 \K_r7_reg[23]  ( .D(K_r6[23]), .CK(n290), .Q(K_r7[23]) );
  DFFQX1 \K_r8_reg[23]  ( .D(K_r7[23]), .CK(n290), .Q(K_r8[23]) );
  DFFQX1 \K_r10_reg[23]  ( .D(K_r9[23]), .CK(n290), .Q(K_r10[23]) );
  DFFQX1 \K_r11_reg[23]  ( .D(K_r10[23]), .CK(n290), .Q(K_r11[23]) );
  DFFQX1 \K_r13_reg[23]  ( .D(K_r12[23]), .CK(n290), .Q(K_r13[23]) );
  DFFQX1 \K_r2_reg[22]  ( .D(K_r1[22]), .CK(n289), .Q(K_r2[22]) );
  DFFQX1 \K_r3_reg[22]  ( .D(K_r2[22]), .CK(n289), .Q(K_r3[22]) );
  DFFQX1 \K_r4_reg[22]  ( .D(K_r3[22]), .CK(n289), .Q(K_r4[22]) );
  DFFQX1 \K_r5_reg[22]  ( .D(K_r4[22]), .CK(n289), .Q(K_r5[22]) );
  DFFQX1 \K_r8_reg[22]  ( .D(K_r7[22]), .CK(n289), .Q(K_r8[22]) );
  DFFQX1 \K_r9_reg[22]  ( .D(K_r8[22]), .CK(n288), .Q(K_r9[22]) );
  DFFQX1 \K_r10_reg[22]  ( .D(K_r9[22]), .CK(n288), .Q(K_r10[22]) );
  DFFQX1 \K_r11_reg[22]  ( .D(K_r10[22]), .CK(n288), .Q(K_r11[22]) );
  DFFQX1 \K_r0_reg[21]  ( .D(K[21]), .CK(n288), .Q(K_r0[21]) );
  DFFQX1 \K_r4_reg[21]  ( .D(K_r3[21]), .CK(n287), .Q(K_r4[21]) );
  DFFQX1 \K_r6_reg[21]  ( .D(K_r5[21]), .CK(n287), .Q(K_r6[21]) );
  DFFQX1 \K_r7_reg[21]  ( .D(K_r6[21]), .CK(n287), .Q(K_r7[21]) );
  DFFQX1 \K_r9_reg[21]  ( .D(K_r8[21]), .CK(n287), .Q(K_r9[21]) );
  DFFQX1 \K_r10_reg[21]  ( .D(K_r9[21]), .CK(n287), .Q(K_r10[21]) );
  DFFQX1 \K_r13_reg[21]  ( .D(K_r12[21]), .CK(n286), .Q(K_r13[21]) );
  DFFQX1 \K_r0_reg[20]  ( .D(K[20]), .CK(n286), .Q(K_r0[20]) );
  DFFQX1 \K_r4_reg[20]  ( .D(K_r3[20]), .CK(n286), .Q(K_r4[20]) );
  DFFQX1 \K_r6_reg[20]  ( .D(K_r5[20]), .CK(n286), .Q(K_r6[20]) );
  DFFQX1 \K_r7_reg[20]  ( .D(K_r6[20]), .CK(n286), .Q(K_r7[20]) );
  DFFQX1 \K_r8_reg[20]  ( .D(K_r7[20]), .CK(n285), .Q(K_r8[20]) );
  DFFQX1 \K_r9_reg[20]  ( .D(K_r8[20]), .CK(n285), .Q(K_r9[20]) );
  DFFQX1 \K_r10_reg[20]  ( .D(K_r9[20]), .CK(n285), .Q(K_r10[20]) );
  DFFQX1 \K_r13_reg[20]  ( .D(K_r12[20]), .CK(n285), .Q(K_r13[20]) );
  DFFQX1 \K_r2_reg[19]  ( .D(K_r1[19]), .CK(n285), .Q(K_r2[19]) );
  DFFQX1 \K_r4_reg[19]  ( .D(K_r3[19]), .CK(n284), .Q(K_r4[19]) );
  DFFQX1 \K_r9_reg[19]  ( .D(K_r8[19]), .CK(n284), .Q(K_r9[19]) );
  DFFQX1 \K_r11_reg[19]  ( .D(K_r10[19]), .CK(n284), .Q(K_r11[19]) );
  DFFQX1 \K_r0_reg[18]  ( .D(K[18]), .CK(n283), .Q(K_r0[18]) );
  DFFQX1 \K_r2_reg[18]  ( .D(K_r1[18]), .CK(n283), .Q(K_r2[18]) );
  DFFQX1 \K_r3_reg[18]  ( .D(K_r2[18]), .CK(n283), .Q(K_r3[18]) );
  DFFQX1 \K_r5_reg[18]  ( .D(K_r4[18]), .CK(n283), .Q(K_r5[18]) );
  DFFQX1 \K_r6_reg[18]  ( .D(K_r5[18]), .CK(n283), .Q(K_r6[18]) );
  DFFQX1 \K_r7_reg[18]  ( .D(K_r6[18]), .CK(n282), .Q(K_r7[18]) );
  DFFQX1 \K_r8_reg[18]  ( .D(K_r7[18]), .CK(n282), .Q(K_r8[18]) );
  DFFQX1 \K_r10_reg[18]  ( .D(K_r9[18]), .CK(n282), .Q(K_r10[18]) );
  DFFQX1 \K_r11_reg[18]  ( .D(K_r10[18]), .CK(n282), .Q(K_r11[18]) );
  DFFQX1 \K_r13_reg[18]  ( .D(K_r12[18]), .CK(n282), .Q(K_r13[18]) );
  DFFQX1 \K_r1_reg[17]  ( .D(K_r0[17]), .CK(n282), .Q(K_r1[17]) );
  DFFQX1 \K_r2_reg[17]  ( .D(K_r1[17]), .CK(n281), .Q(K_r2[17]) );
  DFFQX1 \K_r3_reg[17]  ( .D(K_r2[17]), .CK(n281), .Q(K_r3[17]) );
  DFFQX1 \K_r4_reg[17]  ( .D(K_r3[17]), .CK(n281), .Q(K_r4[17]) );
  DFFQX1 \K_r5_reg[17]  ( .D(K_r4[17]), .CK(n281), .Q(K_r5[17]) );
  DFFQX1 \K_r6_reg[17]  ( .D(K_r5[17]), .CK(n281), .Q(K_r6[17]) );
  DFFQX1 \K_r7_reg[17]  ( .D(K_r6[17]), .CK(n281), .Q(K_r7[17]) );
  DFFQX1 \K_r8_reg[17]  ( .D(K_r7[17]), .CK(n281), .Q(K_r8[17]) );
  DFFQX1 \K_r9_reg[17]  ( .D(K_r8[17]), .CK(n281), .Q(K_r9[17]) );
  DFFQX1 \K_r10_reg[17]  ( .D(K_r9[17]), .CK(n281), .Q(K_r10[17]) );
  DFFQX1 \K_r11_reg[17]  ( .D(K_r10[17]), .CK(n280), .Q(K_r11[17]) );
  DFFQX1 \K_r12_reg[17]  ( .D(K_r11[17]), .CK(n280), .Q(K_r12[17]) );
  DFFQX1 \K_r0_reg[16]  ( .D(K[16]), .CK(n280), .Q(K_r0[16]) );
  DFFQX1 \K_r2_reg[16]  ( .D(K_r1[16]), .CK(n280), .Q(K_r2[16]) );
  DFFQX1 \K_r4_reg[16]  ( .D(K_r3[16]), .CK(n280), .Q(K_r4[16]) );
  DFFQX1 \K_r6_reg[16]  ( .D(K_r5[16]), .CK(n376), .Q(K_r6[16]) );
  DFFQX1 \K_r7_reg[16]  ( .D(K_r6[16]), .CK(clk), .Q(K_r7[16]) );
  DFFQX1 \K_r9_reg[16]  ( .D(K_r8[16]), .CK(clk), .Q(K_r9[16]) );
  DFFQX1 \K_r11_reg[16]  ( .D(K_r10[16]), .CK(n366), .Q(K_r11[16]) );
  DFFQX1 \K_r13_reg[16]  ( .D(K_r12[16]), .CK(n371), .Q(K_r13[16]) );
  DFFQX1 \K_r0_reg[15]  ( .D(K[15]), .CK(n363), .Q(K_r0[15]) );
  DFFQX1 \K_r2_reg[15]  ( .D(K_r1[15]), .CK(n355), .Q(K_r2[15]) );
  DFFQX1 \K_r3_reg[15]  ( .D(K_r2[15]), .CK(n368), .Q(K_r3[15]) );
  DFFQX1 \K_r4_reg[15]  ( .D(K_r3[15]), .CK(n356), .Q(K_r4[15]) );
  DFFQX1 \K_r5_reg[15]  ( .D(K_r4[15]), .CK(n357), .Q(K_r5[15]) );
  DFFQX1 \K_r6_reg[15]  ( .D(K_r5[15]), .CK(n358), .Q(K_r6[15]) );
  DFFQX1 \K_r7_reg[15]  ( .D(K_r6[15]), .CK(n367), .Q(K_r7[15]) );
  DFFQX1 \K_r8_reg[15]  ( .D(K_r7[15]), .CK(n362), .Q(K_r8[15]) );
  DFFQX1 \K_r9_reg[15]  ( .D(K_r8[15]), .CK(n376), .Q(K_r9[15]) );
  DFFQX1 \K_r10_reg[15]  ( .D(K_r9[15]), .CK(n350), .Q(K_r10[15]) );
  DFFQX1 \K_r11_reg[15]  ( .D(K_r10[15]), .CK(n351), .Q(K_r11[15]) );
  DFFQX1 \K_r13_reg[15]  ( .D(K_r12[15]), .CK(n352), .Q(K_r13[15]) );
  DFFQX1 \K_r4_reg[14]  ( .D(K_r3[14]), .CK(n369), .Q(K_r4[14]) );
  DFFQX1 \K_r6_reg[14]  ( .D(K_r5[14]), .CK(n343), .Q(K_r6[14]) );
  DFFQX1 \K_r7_reg[14]  ( .D(K_r6[14]), .CK(n344), .Q(K_r7[14]) );
  DFFQX1 \K_r9_reg[14]  ( .D(K_r8[14]), .CK(n345), .Q(K_r9[14]) );
  DFFQX1 \K_r0_reg[13]  ( .D(K[13]), .CK(n357), .Q(K_r0[13]) );
  DFFQX1 \K_r2_reg[13]  ( .D(K_r1[13]), .CK(n358), .Q(K_r2[13]) );
  DFFQX1 \K_r4_reg[13]  ( .D(K_r3[13]), .CK(n367), .Q(K_r4[13]) );
  DFFQX1 \K_r6_reg[13]  ( .D(K_r5[13]), .CK(n362), .Q(K_r6[13]) );
  DFFQX1 \K_r11_reg[13]  ( .D(K_r10[13]), .CK(n370), .Q(K_r11[13]) );
  DFFQX1 \K_r13_reg[13]  ( .D(K_r12[13]), .CK(n350), .Q(K_r13[13]) );
  DFFQX1 \K_r0_reg[12]  ( .D(K[12]), .CK(n351), .Q(K_r0[12]) );
  DFFQX1 \K_r2_reg[12]  ( .D(K_r1[12]), .CK(n352), .Q(K_r2[12]) );
  DFFQX1 \K_r3_reg[12]  ( .D(K_r2[12]), .CK(n369), .Q(K_r3[12]) );
  DFFQX1 \K_r4_reg[12]  ( .D(K_r3[12]), .CK(n365), .Q(K_r4[12]) );
  DFFQX1 \K_r5_reg[12]  ( .D(K_r4[12]), .CK(n373), .Q(K_r5[12]) );
  DFFQX1 \K_r8_reg[12]  ( .D(K_r7[12]), .CK(n377), .Q(K_r8[12]) );
  DFFQX1 \K_r9_reg[12]  ( .D(K_r8[12]), .CK(n374), .Q(K_r9[12]) );
  DFFQX1 \K_r10_reg[12]  ( .D(K_r9[12]), .CK(n372), .Q(K_r10[12]) );
  DFFQX1 \K_r11_reg[12]  ( .D(K_r10[12]), .CK(n343), .Q(K_r11[12]) );
  DFFQX1 \K_r13_reg[12]  ( .D(K_r12[12]), .CK(n365), .Q(K_r13[12]) );
  DFFQX1 \K_r0_reg[11]  ( .D(K[11]), .CK(n375), .Q(K_r0[11]) );
  DFFQX1 \K_r2_reg[11]  ( .D(K_r1[11]), .CK(n377), .Q(K_r2[11]) );
  DFFQX1 \K_r4_reg[11]  ( .D(K_r3[11]), .CK(n342), .Q(K_r4[11]) );
  DFFQX1 \K_r5_reg[11]  ( .D(K_r4[11]), .CK(n369), .Q(K_r5[11]) );
  DFFQX1 \K_r7_reg[11]  ( .D(K_r6[11]), .CK(n343), .Q(K_r7[11]) );
  DFFQX1 \K_r8_reg[11]  ( .D(K_r7[11]), .CK(n370), .Q(K_r8[11]) );
  DFFQX1 \K_r9_reg[11]  ( .D(K_r8[11]), .CK(n350), .Q(K_r9[11]) );
  DFFQX1 \K_r11_reg[11]  ( .D(K_r10[11]), .CK(n351), .Q(K_r11[11]) );
  DFFQX1 \K_r13_reg[11]  ( .D(K_r12[11]), .CK(n352), .Q(K_r13[11]) );
  DFFQX1 \K_r0_reg[10]  ( .D(K[10]), .CK(n369), .Q(K_r0[10]) );
  DFFQX1 \K_r4_reg[10]  ( .D(K_r3[10]), .CK(n344), .Q(K_r4[10]) );
  DFFQX1 \K_r6_reg[10]  ( .D(K_r5[10]), .CK(n345), .Q(K_r6[10]) );
  DFFQX1 \K_r7_reg[10]  ( .D(K_r6[10]), .CK(n346), .Q(K_r7[10]) );
  DFFQX1 \K_r9_reg[10]  ( .D(K_r8[10]), .CK(n371), .Q(K_r9[10]) );
  DFFQX1 \K_r11_reg[10]  ( .D(K_r10[10]), .CK(n342), .Q(K_r11[10]) );
  DFFQX1 \K_r13_reg[10]  ( .D(K_r12[10]), .CK(n362), .Q(K_r13[10]) );
  DFFQX1 \K_r0_reg[9]  ( .D(K[9]), .CK(n363), .Q(K_r0[9]) );
  DFFQX1 \K_r1_reg[9]  ( .D(K_r0[9]), .CK(n365), .Q(K_r1[9]) );
  DFFQX1 \K_r2_reg[9]  ( .D(K_r1[9]), .CK(clk), .Q(K_r2[9]) );
  DFFQX1 \K_r4_reg[9]  ( .D(K_r3[9]), .CK(n374), .Q(K_r4[9]) );
  DFFQX1 \K_r5_reg[9]  ( .D(K_r4[9]), .CK(n374), .Q(K_r5[9]) );
  DFFQX1 \K_r6_reg[9]  ( .D(K_r5[9]), .CK(n377), .Q(K_r6[9]) );
  DFFQX1 \K_r7_reg[9]  ( .D(K_r6[9]), .CK(n353), .Q(K_r7[9]) );
  DFFQX1 \K_r8_reg[9]  ( .D(K_r7[9]), .CK(n354), .Q(K_r8[9]) );
  DFFQX1 \K_r9_reg[9]  ( .D(K_r8[9]), .CK(n355), .Q(K_r9[9]) );
  DFFQX1 \K_r11_reg[9]  ( .D(K_r10[9]), .CK(n368), .Q(K_r11[9]) );
  DFFQX1 \K_r13_reg[9]  ( .D(K_r12[9]), .CK(n356), .Q(K_r13[9]) );
  DFFQX1 \K_r0_reg[8]  ( .D(K[8]), .CK(n357), .Q(K_r0[8]) );
  DFFQX1 \K_r3_reg[8]  ( .D(K_r2[8]), .CK(n349), .Q(K_r3[8]) );
  DFFQX1 \K_r6_reg[8]  ( .D(K_r5[8]), .CK(n370), .Q(K_r6[8]) );
  DFFQX1 \K_r7_reg[8]  ( .D(K_r6[8]), .CK(n350), .Q(K_r7[8]) );
  DFFQX1 \K_r9_reg[8]  ( .D(K_r8[8]), .CK(n359), .Q(K_r9[8]) );
  DFFQX1 \K_r13_reg[8]  ( .D(K_r12[8]), .CK(n376), .Q(K_r13[8]) );
  DFFQX1 \K_r0_reg[7]  ( .D(K[7]), .CK(n362), .Q(K_r0[7]) );
  DFFQX1 \K_r3_reg[7]  ( .D(K_r2[7]), .CK(n363), .Q(K_r3[7]) );
  DFFQX1 \K_r4_reg[7]  ( .D(K_r3[7]), .CK(n365), .Q(K_r4[7]) );
  DFFQX1 \K_r9_reg[7]  ( .D(K_r8[7]), .CK(n376), .Q(K_r9[7]) );
  DFFQX1 \K_r0_reg[6]  ( .D(K[6]), .CK(n359), .Q(K_r0[6]) );
  DFFQX1 \K_r2_reg[6]  ( .D(K_r1[6]), .CK(n357), .Q(K_r2[6]) );
  DFFQX1 \K_r3_reg[6]  ( .D(K_r2[6]), .CK(n358), .Q(K_r3[6]) );
  DFFQX1 \K_r4_reg[6]  ( .D(K_r3[6]), .CK(n367), .Q(K_r4[6]) );
  DFFQX1 \K_r5_reg[6]  ( .D(K_r4[6]), .CK(n362), .Q(K_r5[6]) );
  DFFQX1 \K_r6_reg[6]  ( .D(K_r5[6]), .CK(n363), .Q(K_r6[6]) );
  DFFQX1 \K_r9_reg[6]  ( .D(K_r8[6]), .CK(n377), .Q(K_r9[6]) );
  DFFQX1 \K_r10_reg[6]  ( .D(K_r9[6]), .CK(n344), .Q(K_r10[6]) );
  DFFQX1 \K_r11_reg[6]  ( .D(K_r10[6]), .CK(n345), .Q(K_r11[6]) );
  DFFQX1 \K_r13_reg[6]  ( .D(K_r12[6]), .CK(n346), .Q(K_r13[6]) );
  DFFQX1 \K_r0_reg[5]  ( .D(K[5]), .CK(n341), .Q(K_r0[5]) );
  DFFQX1 \K_r3_reg[5]  ( .D(K_r2[5]), .CK(n364), .Q(K_r3[5]) );
  DFFQX1 \K_r10_reg[5]  ( .D(K_r9[5]), .CK(n347), .Q(K_r10[5]) );
  DFFQX1 \K_r13_reg[5]  ( .D(K_r12[5]), .CK(n373), .Q(K_r13[5]) );
  DFFQX1 \K_r4_reg[4]  ( .D(K_r3[4]), .CK(n350), .Q(K_r4[4]) );
  DFFQX1 \K_r5_reg[4]  ( .D(K_r4[4]), .CK(n351), .Q(K_r5[4]) );
  DFFQX1 \K_r6_reg[4]  ( .D(K_r5[4]), .CK(n352), .Q(K_r6[4]) );
  DFFQX1 \K_r8_reg[4]  ( .D(K_r7[4]), .CK(n369), .Q(K_r8[4]) );
  DFFQX1 \K_r9_reg[4]  ( .D(K_r8[4]), .CK(n367), .Q(K_r9[4]) );
  DFFQX1 \K_r0_reg[3]  ( .D(K[3]), .CK(n362), .Q(K_r0[3]) );
  DFFQX1 \K_r2_reg[3]  ( .D(K_r1[3]), .CK(n363), .Q(K_r2[3]) );
  DFFQX1 \K_r4_reg[3]  ( .D(K_r3[3]), .CK(n375), .Q(K_r4[3]) );
  DFFQX1 \K_r5_reg[3]  ( .D(K_r4[3]), .CK(n372), .Q(K_r5[3]) );
  DFFQX1 \K_r6_reg[3]  ( .D(K_r5[3]), .CK(n359), .Q(K_r6[3]) );
  DFFQX1 \K_r7_reg[3]  ( .D(K_r6[3]), .CK(n364), .Q(K_r7[3]) );
  DFFQX1 \K_r9_reg[3]  ( .D(K_r8[3]), .CK(n376), .Q(K_r9[3]) );
  DFFQX1 \K_r11_reg[3]  ( .D(K_r10[3]), .CK(n364), .Q(K_r11[3]) );
  DFFQX1 \K_r13_reg[3]  ( .D(K_r12[3]), .CK(n373), .Q(K_r13[3]) );
  DFFQX1 \K_r2_reg[2]  ( .D(K_r1[2]), .CK(n364), .Q(K_r2[2]) );
  DFFQX1 \K_r5_reg[2]  ( .D(K_r4[2]), .CK(n376), .Q(K_r5[2]) );
  DFFQX1 \K_r8_reg[2]  ( .D(K_r7[2]), .CK(n352), .Q(K_r8[2]) );
  DFFQX1 \K_r11_reg[2]  ( .D(K_r10[2]), .CK(n369), .Q(K_r11[2]) );
  DFFQX1 \K_r1_reg[1]  ( .D(K_r0[1]), .CK(n353), .Q(K_r1[1]) );
  DFFQX1 \K_r2_reg[1]  ( .D(K_r1[1]), .CK(n354), .Q(K_r2[1]) );
  DFFQX1 \K_r5_reg[1]  ( .D(K_r4[1]), .CK(n356), .Q(K_r5[1]) );
  DFFQX1 \K_r6_reg[1]  ( .D(K_r5[1]), .CK(n357), .Q(K_r6[1]) );
  DFFQX1 \K_r7_reg[1]  ( .D(K_r6[1]), .CK(n358), .Q(K_r7[1]) );
  DFFQX1 \K_r9_reg[1]  ( .D(K_r8[1]), .CK(n367), .Q(K_r9[1]) );
  DFFQX1 \K_r11_reg[1]  ( .D(K_r10[1]), .CK(n377), .Q(K_r11[1]) );
  DFFQX1 \K_r12_reg[1]  ( .D(K_r11[1]), .CK(n371), .Q(K_r12[1]) );
  DFFQX1 \K_r0_reg[0]  ( .D(K[0]), .CK(n347), .Q(K_r0[0]) );
  DFFQX1 \K_r2_reg[0]  ( .D(K_r1[0]), .CK(n348), .Q(K_r2[0]) );
  DFFQX1 \K_r3_reg[0]  ( .D(K_r2[0]), .CK(n349), .Q(K_r3[0]) );
  DFFQX1 \K_r5_reg[0]  ( .D(K_r4[0]), .CK(n370), .Q(K_r5[0]) );
  DFFQX1 \K_r8_reg[0]  ( .D(K_r7[0]), .CK(n279), .Q(K_r8[0]) );
  DFFQX1 \K_r10_reg[0]  ( .D(K_r9[0]), .CK(n279), .Q(K_r10[0]) );
  DFFQX1 \K_r11_reg[0]  ( .D(K_r10[0]), .CK(n279), .Q(K_r11[0]) );
  DFFQX1 \K_r13_reg[0]  ( .D(K_r12[0]), .CK(n279), .Q(K_r13[0]) );
  DFFQX1 \K_r5_reg[54]  ( .D(K_r4[54]), .CK(n339), .Q(K_r5[54]) );
  DFFQX1 \K_r8_reg[54]  ( .D(K_r7[54]), .CK(n338), .Q(K_r8[54]) );
  DFFQX1 \K_r1_reg[52]  ( .D(K_r0[52]), .CK(n336), .Q(K_r1[52]) );
  DFFQX1 \K_r7_reg[52]  ( .D(K_r6[52]), .CK(n335), .Q(K_r7[52]) );
  DFFQX1 \K_r1_reg[50]  ( .D(K_r0[50]), .CK(n333), .Q(K_r1[50]) );
  DFFQX1 \K_r6_reg[44]  ( .D(K_r5[44]), .CK(n323), .Q(K_r6[44]) );
  DFFQX1 \K_r13_reg[40]  ( .D(K_r12[40]), .CK(n316), .Q(K_r13[40]) );
  DFFQX1 \K_r12_reg[34]  ( .D(K_r11[34]), .CK(n307), .Q(K_r12[34]) );
  DFFQX1 \K_r10_reg[33]  ( .D(K_r9[33]), .CK(n305), .Q(K_r10[33]) );
  DFFQX1 \K_r1_reg[31]  ( .D(K_r0[31]), .CK(n303), .Q(K_r1[31]) );
  DFFQX1 \K_r1_reg[26]  ( .D(K_r0[26]), .CK(n296), .Q(K_r1[26]) );
  DFFQX1 \K_r12_reg[9]  ( .D(K_r11[9]), .CK(n342), .Q(K_r12[9]) );
  DFFQX1 \K_r8_reg[6]  ( .D(K_r7[6]), .CK(n355), .Q(K_r8[6]) );
  DFFQX1 \K_r1_reg[55]  ( .D(K_r0[55]), .CK(n341), .Q(K_r1[55]) );
  DFFQX1 \K_r4_reg[55]  ( .D(K_r3[55]), .CK(n340), .Q(K_r4[55]) );
  DFFQX1 \K_r9_reg[55]  ( .D(K_r8[55]), .CK(n340), .Q(K_r9[55]) );
  DFFQX1 \K_r11_reg[55]  ( .D(K_r10[55]), .CK(n340), .Q(K_r11[55]) );
  DFFQX1 \K_r12_reg[55]  ( .D(K_r11[55]), .CK(n339), .Q(K_r12[55]) );
  DFFQX1 \K_r2_reg[54]  ( .D(K_r1[54]), .CK(n339), .Q(K_r2[54]) );
  DFFQX1 \K_r11_reg[54]  ( .D(K_r10[54]), .CK(n338), .Q(K_r11[54]) );
  DFFQX1 \K_r4_reg[53]  ( .D(K_r3[53]), .CK(n337), .Q(K_r4[53]) );
  DFFQX1 \K_r5_reg[53]  ( .D(K_r4[53]), .CK(n337), .Q(K_r5[53]) );
  DFFQX1 \K_r9_reg[53]  ( .D(K_r8[53]), .CK(n337), .Q(K_r9[53]) );
  DFFQX1 \K_r9_reg[52]  ( .D(K_r8[52]), .CK(n335), .Q(K_r9[52]) );
  DFFQX1 \K_r12_reg[52]  ( .D(K_r11[52]), .CK(n335), .Q(K_r12[52]) );
  DFFQX1 \K_r4_reg[50]  ( .D(K_r3[50]), .CK(n333), .Q(K_r4[50]) );
  DFFQX1 \K_r12_reg[50]  ( .D(K_r11[50]), .CK(n332), .Q(K_r12[50]) );
  DFFQX1 \K_r6_reg[48]  ( .D(K_r5[48]), .CK(n329), .Q(K_r6[48]) );
  DFFQX1 \K_r7_reg[48]  ( .D(K_r6[48]), .CK(n329), .Q(K_r7[48]) );
  DFFQX1 \K_r5_reg[46]  ( .D(K_r4[46]), .CK(n326), .Q(K_r5[46]) );
  DFFQX1 \K_r0_reg[45]  ( .D(K[45]), .CK(n325), .Q(K_r0[45]) );
  DFFQX1 \K_r2_reg[45]  ( .D(K_r1[45]), .CK(n325), .Q(K_r2[45]) );
  DFFQX1 \K_r3_reg[45]  ( .D(K_r2[45]), .CK(n325), .Q(K_r3[45]) );
  DFFQX1 \K_r6_reg[45]  ( .D(K_r5[45]), .CK(n325), .Q(K_r6[45]) );
  DFFQX1 \K_r10_reg[45]  ( .D(K_r9[45]), .CK(n324), .Q(K_r10[45]) );
  DFFQX1 \K_r11_reg[45]  ( .D(K_r10[45]), .CK(n324), .Q(K_r11[45]) );
  DFFQX1 \K_r2_reg[44]  ( .D(K_r1[44]), .CK(n323), .Q(K_r2[44]) );
  DFFQX1 \K_r7_reg[44]  ( .D(K_r6[44]), .CK(n323), .Q(K_r7[44]) );
  DFFQX1 \K_r11_reg[44]  ( .D(K_r10[44]), .CK(n322), .Q(K_r11[44]) );
  DFFQX1 \K_r0_reg[42]  ( .D(K[42]), .CK(n321), .Q(K_r0[42]) );
  DFFQX1 \K_r6_reg[42]  ( .D(K_r5[42]), .CK(n320), .Q(K_r6[42]) );
  DFFQX1 \K_r7_reg[42]  ( .D(K_r6[42]), .CK(n320), .Q(K_r7[42]) );
  DFFQX1 \K_r9_reg[42]  ( .D(K_r8[42]), .CK(n320), .Q(K_r9[42]) );
  DFFQX1 \K_r13_reg[42]  ( .D(K_r12[42]), .CK(n319), .Q(K_r13[42]) );
  DFFQX1 \K_r0_reg[40]  ( .D(K[40]), .CK(n317), .Q(K_r0[40]) );
  DFFQX1 \K_r0_reg[39]  ( .D(K[39]), .CK(n316), .Q(K_r0[39]) );
  DFFQX1 \K_r3_reg[39]  ( .D(K_r2[39]), .CK(n316), .Q(K_r3[39]) );
  DFFQX1 \K_r5_reg[39]  ( .D(K_r4[39]), .CK(n315), .Q(K_r5[39]) );
  DFFQX1 \K_r8_reg[39]  ( .D(K_r7[39]), .CK(n315), .Q(K_r8[39]) );
  DFFQX1 \K_r10_reg[39]  ( .D(K_r9[39]), .CK(n315), .Q(K_r10[39]) );
  DFFQX1 \K_r13_reg[39]  ( .D(K_r12[39]), .CK(n314), .Q(K_r13[39]) );
  DFFQX1 \K_r1_reg[38]  ( .D(K_r0[38]), .CK(n314), .Q(K_r1[38]) );
  DFFQX1 \K_r5_reg[36]  ( .D(K_r4[36]), .CK(n311), .Q(K_r5[36]) );
  DFFQX1 \K_r0_reg[34]  ( .D(K[34]), .CK(n308), .Q(K_r0[34]) );
  DFFQX1 \K_r13_reg[34]  ( .D(K_r12[34]), .CK(n307), .Q(K_r13[34]) );
  DFFQX1 \K_r4_reg[32]  ( .D(K_r3[32]), .CK(n305), .Q(K_r4[32]) );
  DFFQX1 \K_r3_reg[30]  ( .D(K_r2[30]), .CK(n302), .Q(K_r3[30]) );
  DFFQX1 \K_r10_reg[30]  ( .D(K_r9[30]), .CK(n301), .Q(K_r10[30]) );
  DFFQX1 \K_r4_reg[29]  ( .D(K_r3[29]), .CK(n300), .Q(K_r4[29]) );
  DFFQX1 \K_r9_reg[29]  ( .D(K_r8[29]), .CK(n299), .Q(K_r9[29]) );
  DFFQX1 \K_r12_reg[28]  ( .D(K_r11[28]), .CK(n297), .Q(K_r12[28]) );
  DFFQX1 \K_r2_reg[26]  ( .D(K_r1[26]), .CK(n295), .Q(K_r2[26]) );
  DFFQX1 \K_r11_reg[26]  ( .D(K_r10[26]), .CK(n294), .Q(K_r11[26]) );
  DFFQX1 \K_r1_reg[25]  ( .D(K_r0[25]), .CK(n294), .Q(K_r1[25]) );
  DFFQX1 \K_r12_reg[25]  ( .D(K_r11[25]), .CK(n293), .Q(K_r12[25]) );
  DFFQX1 \K_r3_reg[24]  ( .D(K_r2[24]), .CK(n292), .Q(K_r3[24]) );
  DFFQX1 \K_r6_reg[24]  ( .D(K_r5[24]), .CK(n292), .Q(K_r6[24]) );
  DFFQX1 \K_r7_reg[24]  ( .D(K_r6[24]), .CK(n292), .Q(K_r7[24]) );
  DFFQX1 \K_r8_reg[24]  ( .D(K_r7[24]), .CK(n292), .Q(K_r8[24]) );
  DFFQX1 \K_r0_reg[14]  ( .D(K[14]), .CK(n353), .Q(K_r0[14]) );
  DFFQX1 \K_r2_reg[14]  ( .D(K_r1[14]), .CK(n375), .Q(K_r2[14]) );
  DFFQX1 \K_r5_reg[14]  ( .D(K_r4[14]), .CK(n346), .Q(K_r5[14]) );
  DFFQX1 \K_r8_reg[14]  ( .D(K_r7[14]), .CK(n371), .Q(K_r8[14]) );
  DFFQX1 \K_r11_reg[14]  ( .D(K_r10[14]), .CK(n347), .Q(K_r11[14]) );
  DFFQX1 \K_r13_reg[14]  ( .D(K_r12[14]), .CK(n342), .Q(K_r13[14]) );
  DFFQX1 \K_r9_reg[13]  ( .D(K_r8[13]), .CK(n353), .Q(K_r9[13]) );
  DFFQX1 \K_r6_reg[12]  ( .D(K_r5[12]), .CK(n341), .Q(K_r6[12]) );
  DFFQX1 \K_r7_reg[12]  ( .D(K_r6[12]), .CK(n344), .Q(K_r7[12]) );
  DFFQX1 \K_r6_reg[11]  ( .D(K_r5[11]), .CK(n366), .Q(K_r6[11]) );
  DFFQX1 \K_r2_reg[10]  ( .D(K_r1[10]), .CK(n377), .Q(K_r2[10]) );
  DFFQX1 \K_r5_reg[7]  ( .D(K_r4[7]), .CK(n371), .Q(K_r5[7]) );
  DFFQX1 \K_r8_reg[7]  ( .D(K_r7[7]), .CK(n360), .Q(K_r8[7]) );
  DFFQX1 \K_r13_reg[7]  ( .D(K_r12[7]), .CK(n354), .Q(K_r13[7]) );
  DFFQX1 \K_r11_reg[5]  ( .D(K_r10[5]), .CK(n361), .Q(K_r11[5]) );
  DFFQX1 \K_r7_reg[4]  ( .D(K_r6[4]), .CK(n372), .Q(K_r7[4]) );
  DFFQX1 \K_r3_reg[3]  ( .D(K_r2[3]), .CK(n374), .Q(K_r3[3]) );
  DFFQX1 \K_r10_reg[3]  ( .D(K_r9[3]), .CK(n376), .Q(K_r10[3]) );
  DFFQX1 \K_r3_reg[2]  ( .D(K_r2[2]), .CK(n341), .Q(K_r3[2]) );
  DFFQX1 \K_r6_reg[2]  ( .D(K_r5[2]), .CK(n372), .Q(K_r6[2]) );
  DFFQX1 \K_r7_reg[2]  ( .D(K_r6[2]), .CK(n374), .Q(K_r7[2]) );
  DFFQX1 \K_r10_reg[2]  ( .D(K_r9[2]), .CK(n355), .Q(K_r10[2]) );
  DFFQX1 \K_r3_reg[1]  ( .D(K_r2[1]), .CK(n373), .Q(K_r3[1]) );
  DFFQX1 \K_r4_reg[1]  ( .D(K_r3[1]), .CK(n342), .Q(K_r4[1]) );
  DFFQX1 \K_r8_reg[1]  ( .D(K_r7[1]), .CK(n372), .Q(K_r8[1]) );
  DFFQX1 \K_r10_reg[1]  ( .D(K_r9[1]), .CK(n343), .Q(K_r10[1]) );
  DFFQX1 \K_r2_reg[55]  ( .D(K_r1[55]), .CK(n341), .Q(K_r2[55]) );
  DFFQX1 \K_r0_reg[53]  ( .D(K[53]), .CK(n338), .Q(K_r0[53]) );
  DFFQX1 \K_r13_reg[53]  ( .D(K_r12[53]), .CK(n336), .Q(K_r13[53]) );
  DFFQX1 \K_r5_reg[45]  ( .D(K_r4[45]), .CK(n325), .Q(K_r5[45]) );
  DFFQX1 \K_r8_reg[45]  ( .D(K_r7[45]), .CK(n324), .Q(K_r8[45]) );
  DFFQX1 \K_r1_reg[39]  ( .D(K_r0[39]), .CK(n316), .Q(K_r1[39]) );
  DFFQX1 \K_r12_reg[39]  ( .D(K_r11[39]), .CK(n315), .Q(K_r12[39]) );
  DFFQX1 \K_r2_reg[30]  ( .D(K_r1[30]), .CK(n302), .Q(K_r2[30]) );
  DFFQX1 \K_r11_reg[30]  ( .D(K_r10[30]), .CK(n301), .Q(K_r11[30]) );
  DFFQX1 \K_r4_reg[24]  ( .D(K_r3[24]), .CK(n292), .Q(K_r4[24]) );
  DFFQX1 \K_r9_reg[24]  ( .D(K_r8[24]), .CK(n292), .Q(K_r9[24]) );
  DFFQX1 \K_r3_reg[13]  ( .D(K_r2[13]), .CK(n345), .Q(K_r3[13]) );
  DFFQX1 \K_r10_reg[13]  ( .D(K_r9[13]), .CK(n346), .Q(K_r10[13]) );
  DFFQX1 \K_r4_reg[2]  ( .D(K_r3[2]), .CK(n375), .Q(K_r4[2]) );
  DFFQX1 \K_r9_reg[2]  ( .D(K_r8[2]), .CK(n368), .Q(K_r9[2]) );
  DFFQX1 \K_r0_reg[1]  ( .D(K[1]), .CK(n360), .Q(K_r0[1]) );
  DFFQX1 \K_r13_reg[1]  ( .D(K_r12[1]), .CK(n374), .Q(K_r13[1]) );
  BUFX2 U3 ( .A(n240), .Y(n238) );
  CLKBUFX3 U4 ( .A(n358), .Y(n292) );
  CLKBUFX3 U5 ( .A(n355), .Y(n301) );
  CLKBUFX3 U6 ( .A(n355), .Y(n302) );
  CLKBUFX3 U7 ( .A(n350), .Y(n315) );
  CLKBUFX3 U8 ( .A(n350), .Y(n316) );
  CLKBUFX3 U9 ( .A(n347), .Y(n324) );
  CLKBUFX3 U10 ( .A(n347), .Y(n325) );
  CLKBUFX3 U11 ( .A(n343), .Y(n336) );
  CLKBUFX3 U12 ( .A(n343), .Y(n338) );
  CLKBUFX3 U13 ( .A(n375), .Y(n280) );
  CLKBUFX3 U14 ( .A(n373), .Y(n281) );
  CLKBUFX3 U15 ( .A(n361), .Y(n282) );
  CLKBUFX3 U16 ( .A(n361), .Y(n283) );
  CLKBUFX3 U17 ( .A(n361), .Y(n284) );
  CLKBUFX3 U18 ( .A(n360), .Y(n285) );
  CLKBUFX3 U19 ( .A(n360), .Y(n286) );
  CLKBUFX3 U20 ( .A(n360), .Y(n287) );
  CLKBUFX3 U21 ( .A(n359), .Y(n288) );
  CLKBUFX3 U22 ( .A(n359), .Y(n289) );
  CLKBUFX3 U23 ( .A(n359), .Y(n290) );
  CLKBUFX3 U24 ( .A(n358), .Y(n291) );
  CLKBUFX3 U25 ( .A(n358), .Y(n293) );
  CLKBUFX3 U26 ( .A(n357), .Y(n294) );
  CLKBUFX3 U27 ( .A(n357), .Y(n295) );
  CLKBUFX3 U28 ( .A(n357), .Y(n296) );
  CLKBUFX3 U29 ( .A(n356), .Y(n297) );
  CLKBUFX3 U30 ( .A(n356), .Y(n298) );
  CLKBUFX3 U31 ( .A(n356), .Y(n299) );
  CLKBUFX3 U32 ( .A(n355), .Y(n300) );
  CLKBUFX3 U33 ( .A(n354), .Y(n303) );
  CLKBUFX3 U34 ( .A(n354), .Y(n304) );
  CLKBUFX3 U35 ( .A(n354), .Y(n305) );
  CLKBUFX3 U36 ( .A(n353), .Y(n306) );
  CLKBUFX3 U37 ( .A(n353), .Y(n307) );
  CLKBUFX3 U38 ( .A(n353), .Y(n308) );
  CLKBUFX3 U39 ( .A(n352), .Y(n309) );
  CLKBUFX3 U40 ( .A(n352), .Y(n310) );
  CLKBUFX3 U41 ( .A(n352), .Y(n311) );
  CLKBUFX3 U42 ( .A(n351), .Y(n312) );
  CLKBUFX3 U43 ( .A(n351), .Y(n313) );
  CLKBUFX3 U44 ( .A(n351), .Y(n314) );
  CLKBUFX3 U45 ( .A(n350), .Y(n317) );
  CLKBUFX3 U46 ( .A(n349), .Y(n318) );
  CLKBUFX3 U47 ( .A(n349), .Y(n319) );
  CLKBUFX3 U48 ( .A(n349), .Y(n320) );
  CLKBUFX3 U49 ( .A(n348), .Y(n321) );
  CLKBUFX3 U50 ( .A(n348), .Y(n322) );
  CLKBUFX3 U51 ( .A(n348), .Y(n323) );
  CLKBUFX3 U52 ( .A(n347), .Y(n326) );
  CLKBUFX3 U53 ( .A(n346), .Y(n327) );
  CLKBUFX3 U54 ( .A(n346), .Y(n328) );
  CLKBUFX3 U55 ( .A(n346), .Y(n329) );
  CLKBUFX3 U56 ( .A(n345), .Y(n330) );
  CLKBUFX3 U57 ( .A(n345), .Y(n331) );
  CLKBUFX3 U58 ( .A(n345), .Y(n332) );
  CLKBUFX3 U59 ( .A(n344), .Y(n333) );
  CLKBUFX3 U60 ( .A(n344), .Y(n334) );
  CLKBUFX3 U61 ( .A(n344), .Y(n335) );
  CLKBUFX3 U62 ( .A(n343), .Y(n337) );
  CLKBUFX3 U63 ( .A(n342), .Y(n339) );
  CLKBUFX3 U64 ( .A(n342), .Y(n340) );
  CLKBUFX3 U65 ( .A(n342), .Y(n341) );
  CLKBUFX3 U66 ( .A(n363), .Y(n274) );
  CLKBUFX3 U67 ( .A(n363), .Y(n275) );
  CLKBUFX3 U68 ( .A(n363), .Y(n276) );
  CLKBUFX3 U69 ( .A(n362), .Y(n277) );
  CLKBUFX3 U70 ( .A(n362), .Y(n278) );
  CLKBUFX3 U71 ( .A(n362), .Y(n279) );
  CLKBUFX3 U72 ( .A(n366), .Y(n361) );
  CLKBUFX3 U73 ( .A(n366), .Y(n360) );
  CLKBUFX3 U74 ( .A(n366), .Y(n359) );
  CLKBUFX3 U75 ( .A(n367), .Y(n358) );
  CLKBUFX3 U76 ( .A(n367), .Y(n357) );
  CLKBUFX3 U77 ( .A(n367), .Y(n356) );
  CLKBUFX3 U78 ( .A(n368), .Y(n355) );
  CLKBUFX3 U79 ( .A(n368), .Y(n354) );
  CLKBUFX3 U80 ( .A(n368), .Y(n353) );
  CLKBUFX3 U81 ( .A(n369), .Y(n352) );
  CLKBUFX3 U82 ( .A(n369), .Y(n351) );
  CLKBUFX3 U83 ( .A(n369), .Y(n350) );
  CLKBUFX3 U84 ( .A(n370), .Y(n349) );
  CLKBUFX3 U85 ( .A(n370), .Y(n348) );
  CLKBUFX3 U86 ( .A(n370), .Y(n347) );
  CLKBUFX3 U87 ( .A(n371), .Y(n346) );
  CLKBUFX3 U88 ( .A(n371), .Y(n345) );
  CLKBUFX3 U89 ( .A(n371), .Y(n344) );
  CLKBUFX3 U90 ( .A(n372), .Y(n343) );
  CLKBUFX3 U91 ( .A(n372), .Y(n342) );
  CLKBUFX3 U92 ( .A(n364), .Y(n273) );
  CLKBUFX3 U93 ( .A(n365), .Y(n364) );
  CLKBUFX3 U94 ( .A(n341), .Y(n366) );
  CLKBUFX3 U95 ( .A(n375), .Y(n367) );
  CLKBUFX3 U96 ( .A(n375), .Y(n368) );
  CLKBUFX3 U97 ( .A(n374), .Y(n369) );
  CLKBUFX3 U98 ( .A(n374), .Y(n370) );
  CLKBUFX3 U99 ( .A(n373), .Y(n371) );
  CLKBUFX3 U100 ( .A(n365), .Y(n363) );
  CLKBUFX3 U101 ( .A(n365), .Y(n362) );
  CLKBUFX3 U102 ( .A(n373), .Y(n372) );
  CLKBUFX3 U103 ( .A(n377), .Y(n375) );
  CLKBUFX3 U104 ( .A(n377), .Y(n374) );
  CLKBUFX3 U105 ( .A(n377), .Y(n373) );
  CLKBUFX3 U106 ( .A(n376), .Y(n365) );
  CLKBUFX3 U107 ( .A(n375), .Y(n376) );
  CLKBUFX3 U108 ( .A(clk), .Y(n377) );
  CLKINVX1 U109 ( .A(n224), .Y(n8) );
  CLKINVX1 U110 ( .A(n223), .Y(n4) );
  CLKINVX1 U111 ( .A(n223), .Y(n3) );
  CLKINVX1 U112 ( .A(n223), .Y(n6) );
  CLKINVX1 U113 ( .A(n222), .Y(n1) );
  CLKINVX1 U114 ( .A(n223), .Y(n7) );
  CLKINVX1 U115 ( .A(n223), .Y(n5) );
  CLKINVX1 U116 ( .A(n223), .Y(n2) );
  CLKINVX1 U117 ( .A(n224), .Y(n9) );
  CLKINVX1 U118 ( .A(n225), .Y(n16) );
  CLKINVX1 U119 ( .A(n224), .Y(n12) );
  CLKINVX1 U120 ( .A(n224), .Y(n14) );
  CLKINVX1 U121 ( .A(n224), .Y(n10) );
  CLKINVX1 U122 ( .A(n225), .Y(n15) );
  CLKINVX1 U123 ( .A(n224), .Y(n13) );
  CLKINVX1 U124 ( .A(n225), .Y(n17) );
  CLKINVX1 U125 ( .A(n224), .Y(n11) );
  CLKINVX1 U126 ( .A(n225), .Y(n18) );
  CLKINVX1 U127 ( .A(n227), .Y(n33) );
  CLKINVX1 U128 ( .A(n226), .Y(n27) );
  CLKINVX1 U129 ( .A(n227), .Y(n35) );
  CLKINVX1 U130 ( .A(n225), .Y(n20) );
  CLKINVX1 U131 ( .A(n225), .Y(n19) );
  CLKINVX1 U132 ( .A(n226), .Y(n24) );
  CLKINVX1 U133 ( .A(n227), .Y(n32) );
  CLKINVX1 U134 ( .A(n226), .Y(n25) );
  CLKINVX1 U135 ( .A(n226), .Y(n26) );
  CLKINVX1 U136 ( .A(n226), .Y(n28) );
  CLKINVX1 U137 ( .A(n227), .Y(n29) );
  CLKINVX1 U138 ( .A(n226), .Y(n23) );
  CLKINVX1 U139 ( .A(n226), .Y(n22) );
  CLKINVX1 U140 ( .A(n227), .Y(n34) );
  CLKINVX1 U141 ( .A(n225), .Y(n21) );
  CLKINVX1 U142 ( .A(n227), .Y(n31) );
  CLKINVX1 U143 ( .A(n227), .Y(n30) );
  CLKINVX1 U144 ( .A(n231), .Y(n58) );
  CLKINVX1 U145 ( .A(n228), .Y(n38) );
  CLKINVX1 U146 ( .A(n237), .Y(n97) );
  CLKINVX1 U147 ( .A(n228), .Y(n37) );
  CLKINVX1 U148 ( .A(n232), .Y(n60) );
  CLKINVX1 U149 ( .A(n232), .Y(n63) );
  CLKINVX1 U150 ( .A(n230), .Y(n48) );
  CLKINVX1 U151 ( .A(n236), .Y(n93) );
  CLKINVX1 U152 ( .A(n236), .Y(n92) );
  CLKINVX1 U153 ( .A(n236), .Y(n90) );
  CLKINVX1 U154 ( .A(n235), .Y(n85) );
  CLKINVX1 U155 ( .A(n234), .Y(n79) );
  CLKINVX1 U156 ( .A(n234), .Y(n77) );
  CLKINVX1 U157 ( .A(n237), .Y(n98) );
  CLKINVX1 U158 ( .A(n230), .Y(n47) );
  CLKINVX1 U159 ( .A(n231), .Y(n57) );
  CLKINVX1 U160 ( .A(n233), .Y(n68) );
  CLKINVX1 U161 ( .A(n233), .Y(n72) );
  CLKINVX1 U162 ( .A(n230), .Y(n51) );
  CLKINVX1 U163 ( .A(n229), .Y(n39) );
  CLKINVX1 U164 ( .A(n229), .Y(n41) );
  CLKINVX1 U165 ( .A(n237), .Y(n100) );
  CLKINVX1 U166 ( .A(n237), .Y(n94) );
  CLKINVX1 U167 ( .A(n236), .Y(n87) );
  CLKINVX1 U168 ( .A(n235), .Y(n83) );
  CLKINVX1 U169 ( .A(n234), .Y(n74) );
  CLKINVX1 U170 ( .A(n235), .Y(n82) );
  CLKINVX1 U171 ( .A(n234), .Y(n76) );
  CLKINVX1 U172 ( .A(n234), .Y(n78) );
  CLKINVX1 U173 ( .A(n235), .Y(n81) );
  CLKINVX1 U174 ( .A(n228), .Y(n36) );
  CLKINVX1 U175 ( .A(n230), .Y(n49) );
  CLKINVX1 U176 ( .A(n229), .Y(n45) );
  CLKINVX1 U177 ( .A(n232), .Y(n61) );
  CLKINVX1 U178 ( .A(n232), .Y(n64) );
  CLKINVX1 U179 ( .A(n233), .Y(n66) );
  CLKINVX1 U180 ( .A(n233), .Y(n67) );
  CLKINVX1 U181 ( .A(n233), .Y(n70) );
  CLKINVX1 U182 ( .A(n233), .Y(n71) );
  CLKINVX1 U183 ( .A(n233), .Y(n69) );
  CLKINVX1 U184 ( .A(n231), .Y(n55) );
  CLKINVX1 U185 ( .A(n232), .Y(n62) );
  CLKINVX1 U186 ( .A(n232), .Y(n59) );
  CLKINVX1 U187 ( .A(n230), .Y(n52) );
  CLKINVX1 U188 ( .A(n231), .Y(n54) );
  CLKINVX1 U189 ( .A(n229), .Y(n43) );
  CLKINVX1 U190 ( .A(n237), .Y(n99) );
  CLKINVX1 U191 ( .A(n236), .Y(n88) );
  CLKINVX1 U192 ( .A(n235), .Y(n86) );
  CLKINVX1 U193 ( .A(n237), .Y(n96) );
  CLKINVX1 U194 ( .A(n235), .Y(n80) );
  CLKINVX1 U195 ( .A(n235), .Y(n84) );
  CLKINVX1 U196 ( .A(n236), .Y(n89) );
  CLKINVX1 U197 ( .A(n234), .Y(n75) );
  CLKINVX1 U198 ( .A(n236), .Y(n91) );
  CLKINVX1 U199 ( .A(n229), .Y(n40) );
  CLKINVX1 U200 ( .A(n229), .Y(n44) );
  CLKINVX1 U201 ( .A(n234), .Y(n73) );
  CLKINVX1 U202 ( .A(n229), .Y(n42) );
  CLKINVX1 U203 ( .A(n232), .Y(n65) );
  CLKINVX1 U204 ( .A(n230), .Y(n50) );
  CLKINVX1 U205 ( .A(n230), .Y(n46) );
  CLKINVX1 U206 ( .A(n237), .Y(n95) );
  CLKINVX1 U207 ( .A(n231), .Y(n53) );
  CLKINVX1 U208 ( .A(n231), .Y(n56) );
  CLKINVX1 U209 ( .A(n216), .Y(n111) );
  CLKINVX1 U210 ( .A(n217), .Y(n118) );
  CLKINVX1 U211 ( .A(n215), .Y(n103) );
  CLKINVX1 U212 ( .A(n215), .Y(n106) );
  CLKINVX1 U213 ( .A(n215), .Y(n102) );
  CLKINVX1 U214 ( .A(n217), .Y(n116) );
  CLKINVX1 U215 ( .A(n217), .Y(n117) );
  CLKINVX1 U216 ( .A(n215), .Y(n101) );
  CLKINVX1 U217 ( .A(n216), .Y(n110) );
  CLKINVX1 U218 ( .A(n215), .Y(n104) );
  CLKINVX1 U219 ( .A(n216), .Y(n113) );
  CLKINVX1 U220 ( .A(n215), .Y(n105) );
  CLKINVX1 U221 ( .A(n216), .Y(n109) );
  CLKINVX1 U222 ( .A(n217), .Y(n115) );
  CLKINVX1 U223 ( .A(n216), .Y(n108) );
  CLKINVX1 U224 ( .A(n216), .Y(n112) );
  CLKINVX1 U225 ( .A(n216), .Y(n114) );
  CLKINVX1 U226 ( .A(n215), .Y(n107) );
  CLKINVX1 U227 ( .A(n217), .Y(n119) );
  CLKINVX1 U228 ( .A(n221), .Y(n144) );
  CLKINVX1 U229 ( .A(n219), .Y(n132) );
  CLKINVX1 U230 ( .A(n218), .Y(n122) );
  CLKINVX1 U231 ( .A(n219), .Y(n130) );
  CLKINVX1 U232 ( .A(n220), .Y(n141) );
  CLKINVX1 U233 ( .A(n221), .Y(n143) );
  CLKINVX1 U234 ( .A(n221), .Y(n149) );
  CLKINVX1 U235 ( .A(n222), .Y(n154) );
  CLKINVX1 U236 ( .A(n219), .Y(n135) );
  CLKINVX1 U237 ( .A(n221), .Y(n146) );
  CLKINVX1 U238 ( .A(n220), .Y(n137) );
  CLKINVX1 U239 ( .A(n218), .Y(n123) );
  CLKINVX1 U240 ( .A(n217), .Y(n120) );
  CLKINVX1 U241 ( .A(n218), .Y(n126) );
  CLKINVX1 U242 ( .A(n220), .Y(n140) );
  CLKINVX1 U243 ( .A(n221), .Y(n148) );
  CLKINVX1 U244 ( .A(n222), .Y(n153) );
  CLKINVX1 U245 ( .A(n222), .Y(n152) );
  CLKINVX1 U246 ( .A(n219), .Y(n131) );
  CLKINVX1 U247 ( .A(n218), .Y(n128) );
  CLKINVX1 U248 ( .A(n220), .Y(n142) );
  CLKINVX1 U249 ( .A(n223), .Y(n156) );
  CLKINVX1 U250 ( .A(n221), .Y(n145) );
  CLKINVX1 U251 ( .A(n220), .Y(n139) );
  CLKINVX1 U252 ( .A(n218), .Y(n127) );
  CLKINVX1 U253 ( .A(n218), .Y(n124) );
  CLKINVX1 U254 ( .A(n222), .Y(n150) );
  CLKINVX1 U255 ( .A(n221), .Y(n147) );
  CLKINVX1 U256 ( .A(n222), .Y(n151) );
  CLKINVX1 U257 ( .A(n219), .Y(n133) );
  CLKINVX1 U258 ( .A(n220), .Y(n136) );
  CLKINVX1 U259 ( .A(n219), .Y(n129) );
  CLKINVX1 U260 ( .A(n219), .Y(n134) );
  CLKINVX1 U261 ( .A(n218), .Y(n125) );
  CLKINVX1 U262 ( .A(n222), .Y(n155) );
  CLKINVX1 U263 ( .A(n220), .Y(n138) );
  CLKINVX1 U264 ( .A(n217), .Y(n121) );
  CLKBUFX3 U265 ( .A(n248), .Y(n200) );
  CLKBUFX3 U266 ( .A(n253), .Y(n181) );
  CLKBUFX3 U267 ( .A(n255), .Y(n175) );
  CLKBUFX3 U268 ( .A(n249), .Y(n199) );
  CLKBUFX3 U269 ( .A(n252), .Y(n186) );
  CLKBUFX3 U270 ( .A(n254), .Y(n176) );
  CLKBUFX3 U271 ( .A(n250), .Y(n194) );
  CLKBUFX3 U272 ( .A(n251), .Y(n189) );
  CLKBUFX3 U273 ( .A(n255), .Y(n174) );
  CLKBUFX3 U274 ( .A(n251), .Y(n190) );
  CLKBUFX3 U275 ( .A(n251), .Y(n191) );
  CLKBUFX3 U276 ( .A(n249), .Y(n198) );
  CLKBUFX3 U277 ( .A(n248), .Y(n201) );
  CLKBUFX3 U278 ( .A(n248), .Y(n202) );
  CLKBUFX3 U279 ( .A(n256), .Y(n171) );
  CLKBUFX3 U280 ( .A(n251), .Y(n188) );
  CLKBUFX3 U281 ( .A(n252), .Y(n187) );
  CLKBUFX3 U282 ( .A(n253), .Y(n180) );
  CLKBUFX3 U283 ( .A(n254), .Y(n178) );
  CLKBUFX3 U284 ( .A(n255), .Y(n173) );
  CLKBUFX3 U285 ( .A(n248), .Y(n203) );
  CLKBUFX3 U286 ( .A(n254), .Y(n179) );
  CLKBUFX3 U287 ( .A(n252), .Y(n185) );
  CLKBUFX3 U288 ( .A(n256), .Y(n170) );
  CLKBUFX3 U289 ( .A(n250), .Y(n192) );
  CLKBUFX3 U290 ( .A(n250), .Y(n195) );
  CLKBUFX3 U291 ( .A(n250), .Y(n193) );
  CLKBUFX3 U292 ( .A(n249), .Y(n197) );
  CLKBUFX3 U293 ( .A(n249), .Y(n196) );
  CLKBUFX3 U294 ( .A(n253), .Y(n182) );
  CLKBUFX3 U295 ( .A(n256), .Y(n169) );
  CLKBUFX3 U296 ( .A(n253), .Y(n183) );
  CLKBUFX3 U297 ( .A(n252), .Y(n184) );
  CLKBUFX3 U298 ( .A(n255), .Y(n172) );
  CLKBUFX3 U299 ( .A(n254), .Y(n177) );
  CLKBUFX3 U300 ( .A(n246), .Y(n213) );
  CLKBUFX3 U301 ( .A(n246), .Y(n214) );
  CLKBUFX3 U302 ( .A(n169), .Y(n205) );
  CLKBUFX3 U303 ( .A(n226), .Y(n204) );
  CLKBUFX3 U304 ( .A(n239), .Y(n206) );
  CLKBUFX3 U305 ( .A(n247), .Y(n207) );
  CLKBUFX3 U306 ( .A(n247), .Y(n208) );
  CLKBUFX3 U307 ( .A(n247), .Y(n209) );
  CLKBUFX3 U308 ( .A(n246), .Y(n212) );
  CLKBUFX3 U309 ( .A(n247), .Y(n210) );
  CLKBUFX3 U310 ( .A(n246), .Y(n211) );
  CLKBUFX3 U311 ( .A(n258), .Y(n162) );
  CLKBUFX3 U312 ( .A(n257), .Y(n168) );
  CLKBUFX3 U313 ( .A(n258), .Y(n164) );
  CLKBUFX3 U314 ( .A(n257), .Y(n167) );
  CLKBUFX3 U315 ( .A(n257), .Y(n165) );
  CLKBUFX3 U316 ( .A(n258), .Y(n163) );
  CLKBUFX3 U317 ( .A(n257), .Y(n166) );
  CLKBUFX3 U318 ( .A(n259), .Y(n157) );
  CLKBUFX3 U319 ( .A(n259), .Y(n159) );
  CLKBUFX3 U320 ( .A(n259), .Y(n158) );
  CLKBUFX3 U321 ( .A(n259), .Y(n160) );
  CLKBUFX3 U322 ( .A(n258), .Y(n161) );
  CLKBUFX3 U323 ( .A(n239), .Y(n228) );
  CLKBUFX3 U324 ( .A(n241), .Y(n236) );
  CLKBUFX3 U325 ( .A(n241), .Y(n234) );
  CLKBUFX3 U326 ( .A(n238), .Y(n227) );
  CLKBUFX3 U327 ( .A(n242), .Y(n233) );
  CLKBUFX3 U328 ( .A(n243), .Y(n224) );
  CLKBUFX3 U329 ( .A(n244), .Y(n221) );
  CLKBUFX3 U330 ( .A(n241), .Y(n237) );
  CLKBUFX3 U331 ( .A(n244), .Y(n220) );
  CLKBUFX3 U332 ( .A(n243), .Y(n226) );
  CLKBUFX3 U333 ( .A(n242), .Y(n230) );
  CLKBUFX3 U334 ( .A(n239), .Y(n229) );
  CLKBUFX3 U335 ( .A(n244), .Y(n219) );
  CLKBUFX3 U336 ( .A(n245), .Y(n218) );
  CLKBUFX3 U337 ( .A(n242), .Y(n232) );
  CLKBUFX3 U338 ( .A(n245), .Y(n215) );
  CLKBUFX3 U339 ( .A(n242), .Y(n231) );
  CLKBUFX3 U340 ( .A(n245), .Y(n217) );
  CLKBUFX3 U341 ( .A(n243), .Y(n223) );
  CLKBUFX3 U342 ( .A(n241), .Y(n235) );
  CLKBUFX3 U343 ( .A(n244), .Y(n222) );
  CLKBUFX3 U344 ( .A(n243), .Y(n225) );
  CLKBUFX3 U345 ( .A(n245), .Y(n216) );
  CLKBUFX3 U346 ( .A(n263), .Y(n248) );
  CLKBUFX3 U347 ( .A(n262), .Y(n253) );
  CLKBUFX3 U348 ( .A(n261), .Y(n254) );
  CLKBUFX3 U349 ( .A(n262), .Y(n251) );
  CLKBUFX3 U350 ( .A(n261), .Y(n255) );
  CLKBUFX3 U351 ( .A(n263), .Y(n250) );
  CLKBUFX3 U352 ( .A(n263), .Y(n249) );
  CLKBUFX3 U353 ( .A(n237), .Y(n247) );
  CLKBUFX3 U354 ( .A(n261), .Y(n256) );
  CLKBUFX3 U355 ( .A(n262), .Y(n252) );
  CLKBUFX3 U356 ( .A(n235), .Y(n246) );
  CLKBUFX3 U357 ( .A(n240), .Y(n239) );
  CLKBUFX3 U358 ( .A(n265), .Y(n241) );
  CLKBUFX3 U359 ( .A(n260), .Y(n259) );
  CLKBUFX3 U360 ( .A(n264), .Y(n244) );
  CLKBUFX3 U361 ( .A(n265), .Y(n242) );
  CLKBUFX3 U362 ( .A(n264), .Y(n245) );
  CLKBUFX3 U363 ( .A(n260), .Y(n258) );
  CLKBUFX3 U364 ( .A(n264), .Y(n243) );
  CLKBUFX3 U365 ( .A(n260), .Y(n257) );
  CLKBUFX3 U366 ( .A(n268), .Y(n263) );
  CLKBUFX3 U367 ( .A(n268), .Y(n261) );
  CLKBUFX3 U368 ( .A(n268), .Y(n262) );
  CLKBUFX3 U369 ( .A(n266), .Y(n240) );
  CLKBUFX3 U370 ( .A(n267), .Y(n266) );
  CLKBUFX3 U371 ( .A(n270), .Y(n268) );
  CLKBUFX3 U372 ( .A(n267), .Y(n265) );
  CLKBUFX3 U373 ( .A(n267), .Y(n264) );
  CLKBUFX3 U374 ( .A(n269), .Y(n260) );
  CLKBUFX3 U375 ( .A(n270), .Y(n269) );
  CLKBUFX3 U376 ( .A(n272), .Y(n270) );
  CLKBUFX3 U377 ( .A(n271), .Y(n267) );
  CLKBUFX3 U378 ( .A(n272), .Y(n271) );
  OAI22X1 U379 ( .A0(n158), .A1(n427), .B0(n15), .B1(n419), .Y(K14[23]) );
  OAI22X1 U380 ( .A0(n6), .A1(n426), .B0(n163), .B1(n418), .Y(K3[23]) );
  AO22X1 U381 ( .A0(n95), .A1(K_r14[40]), .B0(n257), .B1(K_r14[33]), .Y(
        K16[23]) );
  AO22X1 U382 ( .A0(n206), .A1(K_r13[26]), .B0(n129), .B1(K_r13[47]), .Y(
        K15[23]) );
  AO22X1 U383 ( .A0(n177), .A1(K_r11[55]), .B0(n100), .B1(K_r11[18]), .Y(
        K13[23]) );
  AO22X1 U384 ( .A0(n100), .A1(K_r10[32]), .B0(n267), .B1(K_r10[41]), .Y(
        K12[23]) );
  AO22X1 U385 ( .A0(K_r9[46]), .A1(n28), .B0(K_r9[27]), .B1(n270), .Y(K11[23])
         );
  AO22X1 U386 ( .A0(K_r8[3]), .A1(n35), .B0(K_r8[13]), .B1(n261), .Y(K10[23])
         );
  AO22X1 U387 ( .A0(n193), .A1(K_r7[24]), .B0(n123), .B1(K_r7[17]), .Y(K9[23])
         );
  AO22X1 U388 ( .A0(n26), .A1(K_r6[24]), .B0(n265), .B1(K_r6[17]), .Y(K8[23])
         );
  AO22X1 U389 ( .A0(n237), .A1(K_r5[3]), .B0(K_r5[13]), .B1(n148), .Y(K7[23])
         );
  AO22X1 U390 ( .A0(n238), .A1(K_r4[46]), .B0(K_r4[27]), .B1(n152), .Y(K6[23])
         );
  AO22X1 U391 ( .A0(n219), .A1(K_r3[32]), .B0(n151), .B1(K_r3[41]), .Y(K5[23])
         );
  AO22X1 U392 ( .A0(n72), .A1(K_r2[55]), .B0(n209), .B1(K_r2[18]), .Y(K4[23])
         );
  AO22X1 U393 ( .A0(n59), .A1(K_r0[26]), .B0(n211), .B1(K_r0[47]), .Y(K2[23])
         );
  AO22X1 U394 ( .A0(n187), .A1(K[40]), .B0(n114), .B1(K[33]), .Y(K1[23]) );
  AO22X1 U395 ( .A0(n98), .A1(K_r14[23]), .B0(n209), .B1(K_r14[16]), .Y(
        K16[29]) );
  AO22X1 U396 ( .A0(n40), .A1(K_r13[30]), .B0(n271), .B1(K_r13[9]), .Y(K15[29]) );
  AO22X1 U397 ( .A0(n235), .A1(K_r12[50]), .B0(K_r12[44]), .B1(n145), .Y(
        K14[29]) );
  AO22X1 U398 ( .A0(n176), .A1(K_r11[36]), .B0(n75), .B1(K_r11[31]), .Y(
        K13[29]) );
  AO22X1 U399 ( .A0(n44), .A1(K_r10[45]), .B0(n240), .B1(K_r10[22]), .Y(
        K12[29]) );
  AO22X1 U400 ( .A0(n189), .A1(K_r9[8]), .B0(K_r9[0]), .B1(n124), .Y(K11[29])
         );
  AO22X1 U401 ( .A0(n78), .A1(K_r8[14]), .B0(n213), .B1(K_r8[49]), .Y(K10[29])
         );
  AO22X1 U402 ( .A0(n193), .A1(K_r7[35]), .B0(n127), .B1(K_r7[28]), .Y(K9[29])
         );
  AO22X1 U403 ( .A0(n20), .A1(K_r6[35]), .B0(n211), .B1(K_r6[28]), .Y(K8[29])
         );
  AO22X1 U404 ( .A0(n203), .A1(K_r5[14]), .B0(n120), .B1(K_r5[49]), .Y(K7[29])
         );
  AO22X1 U405 ( .A0(K_r4[8]), .A1(n26), .B0(K_r4[0]), .B1(n269), .Y(K6[29]) );
  AO22X1 U406 ( .A0(n187), .A1(K_r3[45]), .B0(decrypt), .B1(K_r3[22]), .Y(
        K5[29]) );
  AO22X1 U407 ( .A0(n74), .A1(K_r2[36]), .B0(n208), .B1(K_r2[31]), .Y(K4[29])
         );
  AO22X1 U408 ( .A0(K_r1[50]), .A1(n30), .B0(K_r1[44]), .B1(n269), .Y(K3[29])
         );
  AO22X1 U409 ( .A0(n184), .A1(K_r0[30]), .B0(n104), .B1(K_r0[9]), .Y(K2[29])
         );
  AO22X1 U410 ( .A0(n178), .A1(K[23]), .B0(n114), .B1(K[16]), .Y(K1[29]) );
  OAI22X1 U411 ( .A0(n8), .A1(n385), .B0(n166), .B1(n393), .Y(K14[39]) );
  OAI22X1 U412 ( .A0(n162), .A1(n384), .B0(n13), .B1(n392), .Y(K3[39]) );
  AO22X1 U413 ( .A0(K_r14[22]), .A1(n19), .B0(K_r14[15]), .B1(n177), .Y(
        K16[39]) );
  AO22X1 U414 ( .A0(n199), .A1(K_r13[8]), .B0(n116), .B1(K_r13[29]), .Y(
        K15[39]) );
  AO22X1 U415 ( .A0(n175), .A1(K_r11[35]), .B0(n69), .B1(K_r11[2]), .Y(K13[39]) );
  AO22X1 U416 ( .A0(n181), .A1(K_r10[21]), .B0(K_r10[16]), .B1(n137), .Y(
        K12[39]) );
  AO22X1 U417 ( .A0(n92), .A1(K_r9[30]), .B0(n267), .B1(K_r9[7]), .Y(K11[39])
         );
  AO22X1 U418 ( .A0(n81), .A1(K_r8[44]), .B0(n213), .B1(K_r8[52]), .Y(K10[39])
         );
  AO22X1 U419 ( .A0(n191), .A1(K_r7[38]), .B0(K_r7[31]), .B1(n124), .Y(K9[39])
         );
  AO22X1 U420 ( .A0(K_r6[38]), .A1(n24), .B0(K_r6[31]), .B1(n243), .Y(K8[39])
         );
  AO22X1 U421 ( .A0(n202), .A1(K_r5[44]), .B0(n124), .B1(K_r5[52]), .Y(K7[39])
         );
  AO22X1 U422 ( .A0(n241), .A1(K_r4[30]), .B0(n71), .B1(K_r4[7]), .Y(K6[39])
         );
  AO22X1 U423 ( .A0(K_r3[21]), .A1(n26), .B0(K_r3[16]), .B1(n264), .Y(K5[39])
         );
  AO22X1 U424 ( .A0(n72), .A1(K_r2[35]), .B0(n208), .B1(K_r2[2]), .Y(K4[39])
         );
  AO22X1 U425 ( .A0(n61), .A1(K_r0[8]), .B0(n210), .B1(K_r0[29]), .Y(K2[39])
         );
  AO22X1 U426 ( .A0(n176), .A1(K[22]), .B0(K[15]), .B1(n145), .Y(K1[39]) );
  OAI22X1 U427 ( .A0(n160), .A1(n429), .B0(n10), .B1(n421), .Y(K14[11]) );
  OAI22X1 U428 ( .A0(n7), .A1(n428), .B0(n163), .B1(n420), .Y(K3[11]) );
  AO22X1 U429 ( .A0(n194), .A1(K_r14[32]), .B0(K_r14[39]), .B1(n153), .Y(
        K16[11]) );
  AO22X1 U430 ( .A0(K_r13[46]), .A1(n29), .B0(K_r13[25]), .B1(n201), .Y(
        K15[11]) );
  AO22X1 U431 ( .A0(n179), .A1(K_r11[54]), .B0(n77), .B1(K_r11[17]), .Y(
        K13[11]) );
  AO22X1 U432 ( .A0(n185), .A1(K_r10[40]), .B0(n43), .B1(K_r10[6]), .Y(K12[11]) );
  AO22X1 U433 ( .A0(n173), .A1(K_r9[26]), .B0(n74), .B1(K_r9[20]), .Y(K11[11])
         );
  AO22X1 U434 ( .A0(n74), .A1(K_r8[34]), .B0(n254), .B1(K_r8[12]), .Y(K10[11])
         );
  AO22X1 U435 ( .A0(n93), .A1(K_r7[48]), .B0(K_r7[55]), .B1(n245), .Y(K9[11])
         );
  AO22X1 U436 ( .A0(n200), .A1(K_r6[48]), .B0(K_r6[55]), .B1(n140), .Y(K8[11])
         );
  AO22X1 U437 ( .A0(n207), .A1(K_r5[34]), .B0(n19), .B1(K_r5[12]), .Y(K7[11])
         );
  AO22X1 U438 ( .A0(n49), .A1(K_r4[26]), .B0(n205), .B1(K_r4[20]), .Y(K6[11])
         );
  AO22X1 U439 ( .A0(n67), .A1(K_r3[40]), .B0(n164), .B1(K_r3[6]), .Y(K5[11])
         );
  AO22X1 U440 ( .A0(n70), .A1(K_r2[54]), .B0(n209), .B1(K_r2[17]), .Y(K4[11])
         );
  AO22X1 U441 ( .A0(n179), .A1(K_r0[46]), .B0(K_r0[25]), .B1(n141), .Y(K2[11])
         );
  AO22X1 U442 ( .A0(n44), .A1(K[32]), .B0(K[39]), .B1(n189), .Y(K1[11]) );
  AO22X1 U443 ( .A0(n43), .A1(K_r14[13]), .B0(n165), .B1(K_r14[6]), .Y(K16[5])
         );
  AO22X1 U444 ( .A0(n196), .A1(K_r13[24]), .B0(n111), .B1(K_r13[20]), .Y(
        K15[5]) );
  AO22X1 U445 ( .A0(K_r12[34]), .A1(n33), .B0(K_r12[10]), .B1(n202), .Y(K14[5]) );
  AO22X1 U446 ( .A0(n131), .A1(K_r11[48]), .B0(K_r11[53]), .B1(n199), .Y(
        K13[5]) );
  AO22X1 U447 ( .A0(n180), .A1(K_r10[39]), .B0(n28), .B1(K_r10[5]), .Y(K12[5])
         );
  AO22X1 U448 ( .A0(n95), .A1(K_r9[19]), .B0(n255), .B1(K_r9[25]), .Y(K11[5])
         );
  AO22X1 U449 ( .A0(n172), .A1(K_r8[11]), .B0(n35), .B1(K_r8[33]), .Y(K10[5])
         );
  AO22X1 U450 ( .A0(n190), .A1(K_r7[54]), .B0(n39), .B1(K_r7[47]), .Y(K9[5])
         );
  AO22X1 U451 ( .A0(n96), .A1(K_r6[54]), .B0(n253), .B1(K_r6[47]), .Y(K8[5])
         );
  AO22X1 U452 ( .A0(n113), .A1(K_r5[11]), .B0(n260), .B1(K_r5[33]), .Y(K7[5])
         );
  AO22X1 U453 ( .A0(n268), .A1(K_r4[19]), .B0(n36), .B1(K_r4[25]), .Y(K6[5])
         );
  AO22X1 U454 ( .A0(n51), .A1(K_r3[39]), .B0(n205), .B1(K_r3[5]), .Y(K5[5]) );
  AO22X1 U455 ( .A0(n160), .A1(K_r2[48]), .B0(K_r2[53]), .B1(n123), .Y(K4[5])
         );
  AO22X1 U456 ( .A0(n171), .A1(K_r1[34]), .B0(K_r1[10]), .B1(n121), .Y(K3[5])
         );
  AO22X1 U457 ( .A0(n64), .A1(K_r0[24]), .B0(n209), .B1(K_r0[20]), .Y(K2[5])
         );
  AO22X1 U458 ( .A0(n179), .A1(K[13]), .B0(n108), .B1(K[6]), .Y(K1[5]) );
  OAI22X1 U459 ( .A0(n159), .A1(n381), .B0(n13), .B1(n427), .Y(K14[22]) );
  OAI22X1 U460 ( .A0(n7), .A1(n380), .B0(n163), .B1(n426), .Y(K3[22]) );
  AO22X1 U461 ( .A0(n78), .A1(K_r14[32]), .B0(n271), .B1(K_r14[25]), .Y(
        K16[22]) );
  AO22X1 U462 ( .A0(n152), .A1(K_r13[39]), .B0(n269), .B1(K_r13[18]), .Y(
        K15[22]) );
  AO22X1 U463 ( .A0(n30), .A1(K_r11[10]), .B0(K_r11[47]), .B1(n190), .Y(
        K13[22]) );
  AO22X1 U464 ( .A0(n183), .A1(K_r10[33]), .B0(n33), .B1(K_r10[24]), .Y(
        K12[22]) );
  AO22X1 U465 ( .A0(n88), .A1(K_r9[13]), .B0(n262), .B1(K_r9[19]), .Y(K11[22])
         );
  AO22X1 U466 ( .A0(n77), .A1(K_r8[27]), .B0(K_r8[5]), .B1(n244), .Y(K10[22])
         );
  AO22X1 U467 ( .A0(n194), .A1(K_r7[48]), .B0(n126), .B1(K_r7[41]), .Y(K9[22])
         );
  AO22X1 U468 ( .A0(n28), .A1(K_r6[48]), .B0(n270), .B1(K_r6[41]), .Y(K8[22])
         );
  AO22X1 U469 ( .A0(n233), .A1(K_r5[27]), .B0(K_r5[5]), .B1(n149), .Y(K7[22])
         );
  AO22X1 U470 ( .A0(n271), .A1(K_r4[13]), .B0(n94), .B1(K_r4[19]), .Y(K6[22])
         );
  AO22X1 U471 ( .A0(n222), .A1(K_r3[24]), .B0(n155), .B1(K_r3[33]), .Y(K5[22])
         );
  AO22X1 U472 ( .A0(n171), .A1(K_r2[10]), .B0(K_r2[47]), .B1(n129), .Y(K4[22])
         );
  AO22X1 U473 ( .A0(n182), .A1(K_r0[39]), .B0(n105), .B1(K_r0[18]), .Y(K2[22])
         );
  AO22X1 U474 ( .A0(n190), .A1(K[32]), .B0(n116), .B1(K[25]), .Y(K1[22]) );
  OAI22X1 U475 ( .A0(n7), .A1(n423), .B0(n167), .B1(n431), .Y(K14[25]) );
  OAI22X1 U476 ( .A0(n159), .A1(n422), .B0(n11), .B1(n430), .Y(K3[25]) );
  AO22X1 U477 ( .A0(n192), .A1(K_r14[29]), .B0(n109), .B1(K_r14[36]), .Y(
        K16[25]) );
  AO22X1 U478 ( .A0(K_r13[43]), .A1(n27), .B0(K_r13[22]), .B1(n175), .Y(
        K15[25]) );
  AO22X1 U479 ( .A0(n177), .A1(K_r11[49]), .B0(n93), .B1(K_r11[16]), .Y(
        K13[25]) );
  AO22X1 U480 ( .A0(n100), .A1(K_r10[30]), .B0(K_r10[35]), .B1(n264), .Y(
        K12[25]) );
  AO22X1 U481 ( .A0(n189), .A1(K_r9[21]), .B0(n46), .B1(K_r9[44]), .Y(K11[25])
         );
  AO22X1 U482 ( .A0(n170), .A1(K_r8[7]), .B0(n51), .B1(K_r8[31]), .Y(K10[25])
         );
  AO22X1 U483 ( .A0(n193), .A1(K_r7[52]), .B0(n125), .B1(K_r7[45]), .Y(K9[25])
         );
  AO22X1 U484 ( .A0(n198), .A1(K_r6[45]), .B0(n85), .B1(K_r6[52]), .Y(K8[25])
         );
  AO22X1 U485 ( .A0(n105), .A1(K_r5[7]), .B0(n160), .B1(K_r5[31]), .Y(K7[25])
         );
  AO22X1 U486 ( .A0(n44), .A1(K_r4[21]), .B0(n204), .B1(K_r4[44]), .Y(K6[25])
         );
  AO22X1 U487 ( .A0(n218), .A1(K_r3[30]), .B0(K_r3[35]), .B1(n133), .Y(K5[25])
         );
  AO22X1 U488 ( .A0(n73), .A1(K_r2[49]), .B0(n208), .B1(K_r2[16]), .Y(K4[25])
         );
  AO22X1 U489 ( .A0(n183), .A1(K_r0[43]), .B0(K_r0[22]), .B1(n138), .Y(K2[25])
         );
  AO22X1 U490 ( .A0(n48), .A1(K[29]), .B0(n242), .B1(K[36]), .Y(K1[25]) );
  OAI22X1 U491 ( .A0(n159), .A1(n391), .B0(n14), .B1(n409), .Y(K14[33]) );
  OAI22X1 U492 ( .A0(decrypt), .A1(n390), .B0(n164), .B1(n408), .Y(K3[33]) );
  AO22X1 U493 ( .A0(n197), .A1(K_r14[44]), .B0(n114), .B1(K_r14[51]), .Y(
        K16[33]) );
  AO22X1 U494 ( .A0(n201), .A1(K_r13[37]), .B0(K_r13[31]), .B1(n150), .Y(
        K15[33]) );
  AO22X1 U495 ( .A0(n140), .A1(K_r11[0]), .B0(n269), .B1(K_r11[9]), .Y(K13[33]) );
  AO22X1 U496 ( .A0(n182), .A1(K_r10[50]), .B0(K_r10[14]), .B1(n135), .Y(
        K12[33]) );
  AO22X1 U497 ( .A0(n188), .A1(K_r9[36]), .B0(n3), .B1(K_r9[28]), .Y(K11[33])
         );
  AO22X1 U498 ( .A0(n79), .A1(K_r8[42]), .B0(n213), .B1(K_r8[22]), .Y(K10[33])
         );
  AO22X1 U499 ( .A0(n83), .A1(K_r7[1]), .B0(n253), .B1(K_r7[8]), .Y(K9[33]) );
  AO22X1 U500 ( .A0(n197), .A1(K_r6[1]), .B0(n73), .B1(K_r6[8]), .Y(K8[33]) );
  AO22X1 U501 ( .A0(n203), .A1(K_r5[42]), .B0(n89), .B1(K_r5[22]), .Y(K7[33])
         );
  AO22X1 U502 ( .A0(n80), .A1(K_r4[36]), .B0(n204), .B1(K_r4[28]), .Y(K6[33])
         );
  AO22X1 U503 ( .A0(K_r3[50]), .A1(n24), .B0(K_r3[14]), .B1(n160), .Y(K5[33])
         );
  AO22X1 U504 ( .A0(n185), .A1(K_r2[0]), .B0(n41), .B1(K_r2[9]), .Y(K4[33]) );
  AO22X1 U505 ( .A0(K_r0[37]), .A1(n25), .B0(K_r0[31]), .B1(n266), .Y(K2[33])
         );
  AO22X1 U506 ( .A0(n49), .A1(K[44]), .B0(n213), .B1(K[51]), .Y(K1[33]) );
  AO22X1 U507 ( .A0(n41), .A1(K_r14[1]), .B0(K_r14[49]), .B1(n174), .Y(K16[46]) );
  AO22X1 U508 ( .A0(n197), .A1(K_r13[42]), .B0(n110), .B1(K_r13[8]), .Y(
        K15[46]) );
  AO22X1 U509 ( .A0(n198), .A1(K_r12[28]), .B0(K_r12[22]), .B1(n146), .Y(
        K14[46]) );
  AO22X1 U510 ( .A0(n179), .A1(K_r11[14]), .B0(n40), .B1(K_r11[36]), .Y(
        K13[46]) );
  AO22X1 U511 ( .A0(n180), .A1(K_r10[0]), .B0(n27), .B1(K_r10[50]), .Y(K12[46]) );
  AO22X1 U512 ( .A0(n94), .A1(K_r9[9]), .B0(n265), .B1(K_r9[45]), .Y(K11[46])
         );
  AO22X1 U513 ( .A0(n228), .A1(K_r8[31]), .B0(n72), .B1(K_r8[23]), .Y(K10[46])
         );
  AO22X1 U514 ( .A0(n191), .A1(K_r7[44]), .B0(K_r7[37]), .B1(n128), .Y(K9[46])
         );
  AO22X1 U515 ( .A0(K_r6[44]), .A1(n23), .B0(K_r6[37]), .B1(n158), .Y(K8[46])
         );
  AO22X1 U516 ( .A0(n133), .A1(K_r5[31]), .B0(n271), .B1(K_r5[23]), .Y(K7[46])
         );
  AO22X1 U517 ( .A0(n175), .A1(K_r4[9]), .B0(n121), .B1(K_r4[45]), .Y(K6[46])
         );
  AO22X1 U518 ( .A0(n52), .A1(K_r3[0]), .B0(n205), .B1(K_r3[50]), .Y(K5[46])
         );
  AO22X1 U519 ( .A0(n69), .A1(K_r2[14]), .B0(n207), .B1(K_r2[36]), .Y(K4[46])
         );
  AO22X1 U520 ( .A0(K_r1[28]), .A1(n34), .B0(K_r1[22]), .B1(n256), .Y(K3[46])
         );
  AO22X1 U521 ( .A0(n63), .A1(K_r0[42]), .B0(n209), .B1(K_r0[8]), .Y(K2[46])
         );
  AO22X1 U522 ( .A0(n178), .A1(K[1]), .B0(K[49]), .B1(n142), .Y(K1[46]) );
  AO22X1 U523 ( .A0(n201), .A1(K_r14[36]), .B0(K_r14[43]), .B1(n155), .Y(
        K16[44]) );
  AO22X1 U524 ( .A0(n198), .A1(K_r13[29]), .B0(n117), .B1(K_r13[50]), .Y(
        K15[44]) );
  AO22X1 U525 ( .A0(K_r12[9]), .A1(n30), .B0(K_r12[15]), .B1(n198), .Y(K14[44]) );
  AO22X1 U526 ( .A0(n141), .A1(K_r11[23]), .B0(n270), .B1(K_r11[1]), .Y(
        K13[44]) );
  AO22X1 U527 ( .A0(n23), .A1(K_r10[37]), .B0(n262), .B1(K_r10[42]), .Y(
        K12[44]) );
  AO22X1 U528 ( .A0(n187), .A1(K_r9[28]), .B0(n103), .B1(K_r9[51]), .Y(K11[44]) );
  AO22X1 U529 ( .A0(n228), .A1(K_r8[14]), .B0(n99), .B1(K_r8[38]), .Y(K10[44])
         );
  AO22X1 U530 ( .A0(K_r7[52]), .A1(n31), .B0(K_r7[0]), .B1(n264), .Y(K9[44])
         );
  AO22X1 U531 ( .A0(n196), .A1(K_r6[52]), .B0(K_r6[0]), .B1(n132), .Y(K8[44])
         );
  AO22X1 U532 ( .A0(n148), .A1(K_r5[14]), .B0(n168), .B1(K_r5[38]), .Y(K7[44])
         );
  AO22X1 U533 ( .A0(n38), .A1(K_r4[28]), .B0(n166), .B1(K_r4[51]), .Y(K6[44])
         );
  AO22X1 U534 ( .A0(n222), .A1(K_r3[37]), .B0(n99), .B1(K_r3[42]), .Y(K5[44])
         );
  AO22X1 U535 ( .A0(n161), .A1(K_r2[23]), .B0(n21), .B1(K_r2[1]), .Y(K4[44])
         );
  AO22X1 U536 ( .A0(n163), .A1(K_r1[9]), .B0(K_r1[15]), .B1(n123), .Y(K3[44])
         );
  AO22X1 U537 ( .A0(n62), .A1(K_r0[29]), .B0(n210), .B1(K_r0[50]), .Y(K2[44])
         );
  AO22X1 U538 ( .A0(n52), .A1(K[36]), .B0(K[43]), .B1(n191), .Y(K1[44]) );
  AO22X1 U539 ( .A0(n91), .A1(K_r14[14]), .B0(n166), .B1(K_r14[7]), .Y(K16[31]) );
  AO22X1 U540 ( .A0(n100), .A1(K_r13[21]), .B0(n240), .B1(K_r13[0]), .Y(
        K15[31]) );
  OAI22X1 U541 ( .A0(n3), .A1(n391), .B0(n165), .B1(n399), .Y(K14[31]) );
  AO22X1 U542 ( .A0(n176), .A1(K_r11[31]), .B0(n149), .B1(K_r11[49]), .Y(
        K13[31]) );
  AO22X1 U543 ( .A0(K_r10[8]), .A1(n21), .B0(K_r10[44]), .B1(n256), .Y(K12[31]) );
  AO22X1 U544 ( .A0(n90), .A1(K_r9[22]), .B0(n181), .B1(K_r9[30]), .Y(K11[31])
         );
  AO22X1 U545 ( .A0(K_r8[36]), .A1(n30), .B0(K_r8[16]), .B1(n254), .Y(K10[31])
         );
  AO22X1 U546 ( .A0(n192), .A1(K_r7[2]), .B0(n146), .B1(K_r7[50]), .Y(K9[31])
         );
  AO22X1 U547 ( .A0(n19), .A1(K_r6[2]), .B0(n201), .B1(K_r6[50]), .Y(K8[31])
         );
  AO22X1 U548 ( .A0(n203), .A1(K_r5[36]), .B0(K_r5[16]), .B1(n147), .Y(K7[31])
         );
  AO22X1 U549 ( .A0(n181), .A1(K_r4[22]), .B0(n129), .B1(K_r4[30]), .Y(K6[31])
         );
  AO22X1 U550 ( .A0(n197), .A1(K_r3[8]), .B0(K_r3[44]), .B1(n136), .Y(K5[31])
         );
  AO22X1 U551 ( .A0(n42), .A1(K_r2[31]), .B0(n208), .B1(K_r2[49]), .Y(K4[31])
         );
  OAI22X1 U552 ( .A0(n157), .A1(n390), .B0(n12), .B1(n398), .Y(K3[31]) );
  AO22X1 U553 ( .A0(n185), .A1(K_r0[21]), .B0(n102), .B1(K_r0[0]), .Y(K2[31])
         );
  AO22X1 U554 ( .A0(n175), .A1(K[14]), .B0(n112), .B1(K[7]), .Y(K1[31]) );
  AO22X1 U555 ( .A0(n191), .A1(K_r14[54]), .B0(n105), .B1(K_r14[4]), .Y(
        K16[19]) );
  AO22X1 U556 ( .A0(n262), .A1(K_r13[47]), .B0(n24), .B1(K_r13[11]), .Y(
        K15[19]) );
  AO22X1 U557 ( .A0(n135), .A1(K_r12[25]), .B0(K_r12[33]), .B1(n271), .Y(
        K14[19]) );
  AO22X1 U558 ( .A0(n27), .A1(K_r11[39]), .B0(n261), .B1(K_r11[19]), .Y(
        K13[19]) );
  AO22X1 U559 ( .A0(n184), .A1(K_r10[5]), .B0(n35), .B1(K_r10[53]), .Y(K12[19]) );
  AO22X1 U560 ( .A0(n87), .A1(K_r9[10]), .B0(K_r9[48]), .B1(n259), .Y(K11[19])
         );
  AO22X1 U561 ( .A0(n76), .A1(K_r8[24]), .B0(n260), .B1(K_r8[34]), .Y(K10[19])
         );
  AO22X1 U562 ( .A0(K_r7[13]), .A1(n29), .B0(n260), .B1(K_r7[20]), .Y(K9[19])
         );
  AO22X1 U563 ( .A0(n199), .A1(K_r6[13]), .B0(n97), .B1(K_r6[20]), .Y(K8[19])
         );
  AO22X1 U564 ( .A0(n256), .A1(K_r5[24]), .B0(n145), .B1(K_r5[34]), .Y(K7[19])
         );
  AO22X1 U565 ( .A0(n202), .A1(K_r4[10]), .B0(K_r4[48]), .B1(n150), .Y(K6[19])
         );
  AO22X1 U566 ( .A0(n64), .A1(K_r3[5]), .B0(n163), .B1(K_r3[53]), .Y(K5[19])
         );
  AO22X1 U567 ( .A0(n240), .A1(K_r2[39]), .B0(n119), .B1(K_r2[19]), .Y(K4[19])
         );
  AO22X1 U568 ( .A0(n256), .A1(K_r1[25]), .B0(K_r1[33]), .B1(n127), .Y(K3[19])
         );
  AO22X1 U569 ( .A0(n57), .A1(K_r0[47]), .B0(n211), .B1(K_r0[11]), .Y(K2[19])
         );
  AO22X1 U570 ( .A0(n46), .A1(K[54]), .B0(n239), .B1(K[4]), .Y(K1[19]) );
  AO22X1 U571 ( .A0(n197), .A1(K_r14[28]), .B0(n68), .B1(K_r14[35]), .Y(
        K16[35]) );
  AO22X1 U572 ( .A0(n67), .A1(K_r13[42]), .B0(n272), .B1(K_r13[21]), .Y(
        K15[35]) );
  AO22X1 U573 ( .A0(n138), .A1(K_r12[1]), .B0(K_r12[7]), .B1(n197), .Y(K14[35]) );
  AO22X1 U574 ( .A0(n175), .A1(K_r11[52]), .B0(n5), .B1(K_r11[15]), .Y(K13[35]) );
  AO22X1 U575 ( .A0(n182), .A1(K_r10[38]), .B0(n11), .B1(K_r10[29]), .Y(
        K12[35]) );
  AO22X1 U576 ( .A0(n188), .A1(K_r9[51]), .B0(n6), .B1(K_r9[43]), .Y(K11[35])
         );
  AO22X1 U577 ( .A0(n80), .A1(K_r8[2]), .B0(K_r8[37]), .B1(n258), .Y(K10[35])
         );
  AO22X1 U578 ( .A0(n83), .A1(K_r7[16]), .B0(n176), .B1(K_r7[23]), .Y(K9[35])
         );
  AO22X1 U579 ( .A0(n197), .A1(K_r6[16]), .B0(n119), .B1(K_r6[23]), .Y(K8[35])
         );
  AO22X1 U580 ( .A0(n202), .A1(K_r5[2]), .B0(K_r5[37]), .B1(n145), .Y(K7[35])
         );
  AO22X1 U581 ( .A0(n79), .A1(K_r4[51]), .B0(n204), .B1(K_r4[43]), .Y(K6[35])
         );
  AO22X1 U582 ( .A0(n58), .A1(K_r3[38]), .B0(n206), .B1(K_r3[29]), .Y(K5[35])
         );
  AO22X1 U583 ( .A0(n73), .A1(K_r2[52]), .B0(n208), .B1(K_r2[15]), .Y(K4[35])
         );
  AO22X1 U584 ( .A0(n169), .A1(K_r1[1]), .B0(K_r1[7]), .B1(n120), .Y(K3[35])
         );
  AO22X1 U585 ( .A0(n186), .A1(K_r0[42]), .B0(n102), .B1(K_r0[21]), .Y(K2[35])
         );
  AO22X1 U586 ( .A0(n50), .A1(K[28]), .B0(n212), .B1(K[35]), .Y(K1[35]) );
  AO22X1 U587 ( .A0(K_r14[52]), .A1(n27), .B0(K_r14[45]), .B1(n244), .Y(
        K16[30]) );
  AO22X1 U588 ( .A0(n77), .A1(K_r13[0]), .B0(n259), .B1(K_r13[38]), .Y(K15[30]) );
  OAI22X1 U589 ( .A0(n8), .A1(n383), .B0(n167), .B1(n415), .Y(K14[30]) );
  AO22X1 U590 ( .A0(n176), .A1(K_r11[37]), .B0(K_r11[28]), .B1(n141), .Y(
        K13[30]) );
  AO22X1 U591 ( .A0(n45), .A1(K_r10[42]), .B0(n183), .B1(K_r10[23]), .Y(
        K12[30]) );
  AO22X1 U592 ( .A0(n90), .A1(K_r9[1]), .B0(n182), .B1(K_r9[9]), .Y(K11[30])
         );
  AO22X1 U593 ( .A0(n170), .A1(K_r8[50]), .B0(n86), .B1(K_r8[15]), .Y(K10[30])
         );
  AO22X1 U594 ( .A0(n193), .A1(K_r7[36]), .B0(K_r7[29]), .B1(n119), .Y(K9[30])
         );
  AO22X1 U595 ( .A0(K_r6[36]), .A1(n20), .B0(K_r6[29]), .B1(n161), .Y(K8[30])
         );
  AO22X1 U596 ( .A0(n117), .A1(K_r5[50]), .B0(n226), .B1(K_r5[15]), .Y(K7[30])
         );
  AO22X1 U597 ( .A0(n170), .A1(K_r4[1]), .B0(n53), .B1(K_r4[9]), .Y(K6[30]) );
  AO22X1 U598 ( .A0(n196), .A1(K_r3[42]), .B0(decrypt), .B1(K_r3[23]), .Y(
        K5[30]) );
  AO22X1 U599 ( .A0(K_r2[37]), .A1(n92), .B0(K_r2[28]), .B1(n229), .Y(K4[30])
         );
  OAI22X1 U600 ( .A0(n157), .A1(n382), .B0(n15), .B1(n414), .Y(K3[30]) );
  AO22X1 U601 ( .A0(n184), .A1(K_r0[0]), .B0(n102), .B1(K_r0[38]), .Y(K2[30])
         );
  AO22X1 U602 ( .A0(n176), .A1(K[52]), .B0(K[45]), .B1(n149), .Y(K1[30]) );
  AO22X1 U603 ( .A0(K_r14[17]), .A1(n24), .B0(K_r14[10]), .B1(n158), .Y(
        K16[17]) );
  AO22X1 U604 ( .A0(n174), .A1(K_r13[3]), .B0(n25), .B1(K_r13[24]), .Y(K15[17]) );
  OAI22X1 U605 ( .A0(n5), .A1(n389), .B0(n165), .B1(n417), .Y(K14[17]) );
  AO22X1 U606 ( .A0(n178), .A1(K_r11[32]), .B0(K_r11[27]), .B1(n138), .Y(
        K13[17]) );
  AO22X1 U607 ( .A0(n98), .A1(K_r10[41]), .B0(n256), .B1(K_r10[18]), .Y(
        K12[17]) );
  AO22X1 U608 ( .A0(n87), .A1(K_r9[55]), .B0(n268), .B1(K_r9[4]), .Y(K11[17])
         );
  AO22X1 U609 ( .A0(n76), .A1(K_r8[12]), .B0(n269), .B1(K_r8[47]), .Y(K10[17])
         );
  AO22X1 U610 ( .A0(n194), .A1(K_r7[33]), .B0(K_r7[26]), .B1(n121), .Y(K9[17])
         );
  AO22X1 U611 ( .A0(K_r6[33]), .A1(n27), .B0(K_r6[26]), .B1(n261), .Y(K8[17])
         );
  AO22X1 U612 ( .A0(n240), .A1(K_r5[12]), .B0(n23), .B1(K_r5[47]), .Y(K7[17])
         );
  AO22X1 U613 ( .A0(n203), .A1(K_r4[55]), .B0(n83), .B1(K_r4[4]), .Y(K6[17])
         );
  AO22X1 U614 ( .A0(n239), .A1(K_r3[41]), .B0(n153), .B1(K_r3[18]), .Y(K5[17])
         );
  AO22X1 U615 ( .A0(K_r2[32]), .A1(n35), .B0(K_r2[27]), .B1(n257), .Y(K4[17])
         );
  OAI22X1 U616 ( .A0(n158), .A1(n388), .B0(n14), .B1(n416), .Y(K3[17]) );
  AO22X1 U617 ( .A0(n56), .A1(K_r0[3]), .B0(n211), .B1(K_r0[24]), .Y(K2[17])
         );
  AO22X1 U618 ( .A0(n215), .A1(K[17]), .B0(K[10]), .B1(n151), .Y(K1[17]) );
  AO22X1 U619 ( .A0(n191), .A1(K_r14[40]), .B0(n107), .B1(K_r14[47]), .Y(
        K16[1]) );
  AO22X1 U620 ( .A0(n107), .A1(K_r13[54]), .B0(n178), .B1(K_r13[33]), .Y(
        K15[1]) );
  OAI22X1 U621 ( .A0(n5), .A1(n413), .B0(n162), .B1(n421), .Y(K14[1]) );
  AO22X1 U622 ( .A0(n178), .A1(K_r11[5]), .B0(K_r11[25]), .B1(n139), .Y(K13[1]) );
  AO22X1 U623 ( .A0(n99), .A1(K_r10[39]), .B0(n253), .B1(K_r10[48]), .Y(K12[1]) );
  AO22X1 U624 ( .A0(n88), .A1(K_r9[53]), .B0(n263), .B1(K_r9[34]), .Y(K11[1])
         );
  AO22X1 U625 ( .A0(n169), .A1(K_r8[20]), .B0(K_r8[10]), .B1(n133), .Y(K10[1])
         );
  AO22X1 U626 ( .A0(n89), .A1(K_r7[24]), .B0(n228), .B1(K_r7[6]), .Y(K9[1]) );
  AO22X1 U627 ( .A0(n199), .A1(K_r6[24]), .B0(n58), .B1(K_r6[6]), .Y(K8[1]) );
  AO22X1 U628 ( .A0(K_r5[20]), .A1(n29), .B0(K_r5[10]), .B1(n267), .Y(K7[1])
         );
  AO22X1 U629 ( .A0(n169), .A1(K_r4[53]), .B0(n57), .B1(K_r4[34]), .Y(K6[1])
         );
  AO22X1 U630 ( .A0(n239), .A1(K_r3[39]), .B0(n64), .B1(K_r3[48]), .Y(K5[1])
         );
  AO22X1 U631 ( .A0(K_r2[5]), .A1(n32), .B0(K_r2[25]), .B1(n210), .Y(K4[1]) );
  OAI22X1 U632 ( .A0(n158), .A1(n412), .B0(n17), .B1(n420), .Y(K3[1]) );
  AO22X1 U633 ( .A0(n182), .A1(K_r0[54]), .B0(n106), .B1(K_r0[33]), .Y(K2[1])
         );
  AO22X1 U634 ( .A0(n46), .A1(K[40]), .B0(n248), .B1(K[47]), .Y(K1[1]) );
  AO22X1 U635 ( .A0(n190), .A1(K_r14[48]), .B0(n108), .B1(K_r14[55]), .Y(
        K16[20]) );
  AO22X1 U636 ( .A0(n271), .A1(K_r13[41]), .B0(n9), .B1(K_r13[5]), .Y(K15[20])
         );
  OAI22X1 U637 ( .A0(n6), .A1(n405), .B0(n166), .B1(n413), .Y(K14[20]) );
  AO22X1 U638 ( .A0(n177), .A1(K_r11[13]), .B0(K_r11[33]), .B1(n139), .Y(
        K13[20]) );
  AO22X1 U639 ( .A0(n184), .A1(K_r10[24]), .B0(K_r10[47]), .B1(n135), .Y(
        K12[20]) );
  AO22X1 U640 ( .A0(n88), .A1(K_r9[4]), .B0(n250), .B1(K_r9[10]), .Y(K11[20])
         );
  AO22X1 U641 ( .A0(n167), .A1(K_r8[53]), .B0(n49), .B1(K_r8[18]), .Y(K10[20])
         );
  AO22X1 U642 ( .A0(n89), .A1(K_r7[32]), .B0(n247), .B1(K_r7[39]), .Y(K9[20])
         );
  AO22X1 U643 ( .A0(n199), .A1(K_r6[32]), .B0(n92), .B1(K_r6[39]), .Y(K8[20])
         );
  AO22X1 U644 ( .A0(n24), .A1(K_r5[53]), .B0(n220), .B1(K_r5[18]), .Y(K7[20])
         );
  AO22X1 U645 ( .A0(n168), .A1(K_r4[4]), .B0(n96), .B1(K_r4[10]), .Y(K6[20])
         );
  AO22X1 U646 ( .A0(n63), .A1(K_r3[24]), .B0(K_r3[47]), .B1(n251), .Y(K5[20])
         );
  AO22X1 U647 ( .A0(n71), .A1(K_r2[13]), .B0(K_r2[33]), .B1(n253), .Y(K4[20])
         );
  OAI22X1 U648 ( .A0(n158), .A1(n404), .B0(n17), .B1(n412), .Y(K3[20]) );
  AO22X1 U649 ( .A0(n58), .A1(K_r0[41]), .B0(n211), .B1(K_r0[5]), .Y(K2[20])
         );
  AO22X1 U650 ( .A0(n47), .A1(K[48]), .B0(n268), .B1(K[55]), .Y(K1[20]) );
  AO22X1 U651 ( .A0(n43), .A1(K_r14[6]), .B0(n254), .B1(K_r14[24]), .Y(K16[8])
         );
  AO22X1 U652 ( .A0(n46), .A1(K_r13[13]), .B0(K_r13[17]), .B1(n253), .Y(K15[8]) );
  OAI22X1 U653 ( .A0(n2), .A1(n429), .B0(n163), .B1(n405), .Y(K14[8]) );
  AO22X1 U654 ( .A0(n182), .A1(K_r11[46]), .B0(n44), .B1(K_r11[41]), .Y(K13[8]) );
  AO22X1 U655 ( .A0(n48), .A1(K_r10[55]), .B0(n270), .B1(K_r10[32]), .Y(K12[8]) );
  AO22X1 U656 ( .A0(n96), .A1(K_r9[12]), .B0(K_r9[18]), .B1(n245), .Y(K11[8])
         );
  AO22X1 U657 ( .A0(n173), .A1(K_r8[4]), .B0(n155), .B1(K_r8[26]), .Y(K10[8])
         );
  AO22X1 U658 ( .A0(n174), .A1(K_r7[47]), .B0(n145), .B1(K_r7[40]), .Y(K9[8])
         );
  AO22X1 U659 ( .A0(n94), .A1(K_r6[47]), .B0(n210), .B1(K_r6[40]), .Y(K8[8])
         );
  AO22X1 U660 ( .A0(n114), .A1(K_r5[4]), .B0(n166), .B1(K_r5[26]), .Y(K7[8])
         );
  AO22X1 U661 ( .A0(n173), .A1(K_r4[12]), .B0(K_r4[18]), .B1(n151), .Y(K6[8])
         );
  AO22X1 U662 ( .A0(n247), .A1(K_r3[55]), .B0(n82), .B1(K_r3[32]), .Y(K5[8])
         );
  AO22X1 U663 ( .A0(n68), .A1(K_r2[46]), .B0(n207), .B1(K_r2[41]), .Y(K4[8])
         );
  OAI22X1 U664 ( .A0(n161), .A1(n428), .B0(n10), .B1(n404), .Y(K3[8]) );
  AO22X1 U665 ( .A0(n174), .A1(K_r0[13]), .B0(K_r0[17]), .B1(n125), .Y(K2[8])
         );
  AO22X1 U666 ( .A0(n179), .A1(K[6]), .B0(n107), .B1(K[24]), .Y(K1[8]) );
  AO22X1 U667 ( .A0(n194), .A1(K_r14[14]), .B0(n61), .B1(K_r14[21]), .Y(
        K16[27]) );
  AO22X1 U668 ( .A0(n230), .A1(K_r13[7]), .B0(n50), .B1(K_r13[28]), .Y(K15[27]) );
  AO22X1 U669 ( .A0(n174), .A1(K_r12[52]), .B0(K_r12[42]), .B1(n144), .Y(
        K14[27]) );
  AO22X1 U670 ( .A0(n102), .A1(K_r11[1]), .B0(n270), .B1(K_r11[38]), .Y(
        K13[27]) );
  AO22X1 U671 ( .A0(n183), .A1(K_r10[51]), .B0(n12), .B1(K_r10[15]), .Y(
        K12[27]) );
  AO22X1 U672 ( .A0(n89), .A1(K_r9[29]), .B0(n231), .B1(K_r9[37]), .Y(K11[27])
         );
  AO22X1 U673 ( .A0(n169), .A1(K_r8[23]), .B0(K_r8[43]), .B1(n130), .Y(K10[27]) );
  AO22X1 U674 ( .A0(n85), .A1(K_r7[2]), .B0(n246), .B1(K_r7[9]), .Y(K9[27]) );
  AO22X1 U675 ( .A0(n198), .A1(K_r6[2]), .B0(n14), .B1(K_r6[9]), .Y(K8[27]) );
  AO22X1 U676 ( .A0(n156), .A1(K_r5[23]), .B0(K_r5[43]), .B1(n265), .Y(K7[27])
         );
  AO22X1 U677 ( .A0(n186), .A1(K_r4[29]), .B0(n16), .B1(K_r4[37]), .Y(K6[27])
         );
  AO22X1 U678 ( .A0(n60), .A1(K_r3[51]), .B0(n206), .B1(K_r3[15]), .Y(K5[27])
         );
  AO22X1 U679 ( .A0(n173), .A1(K_r2[1]), .B0(n118), .B1(K_r2[38]), .Y(K4[27])
         );
  AO22X1 U680 ( .A0(K_r1[52]), .A1(n32), .B0(K_r1[42]), .B1(n248), .Y(K3[27])
         );
  AO22X1 U681 ( .A0(n59), .A1(K_r0[7]), .B0(n211), .B1(K_r0[28]), .Y(K2[27])
         );
  AO22X1 U682 ( .A0(n48), .A1(K[14]), .B0(n255), .B1(K[21]), .Y(K1[27]) );
  AO22X1 U683 ( .A0(n200), .A1(K_r14[31]), .B0(K_r14[38]), .B1(n156), .Y(
        K16[42]) );
  AO22X1 U684 ( .A0(n36), .A1(K_r13[45]), .B0(n242), .B1(K_r13[51]), .Y(
        K15[42]) );
  AO22X1 U685 ( .A0(n131), .A1(K_r11[14]), .B0(n238), .B1(K_r11[23]), .Y(
        K13[42]) );
  AO22X1 U686 ( .A0(n57), .A1(K_r10[28]), .B0(K_r10[9]), .B1(n252), .Y(K12[42]) );
  AO22X1 U687 ( .A0(n93), .A1(K_r9[42]), .B0(n266), .B1(K_r9[50]), .Y(K11[42])
         );
  AO22X1 U688 ( .A0(n82), .A1(K_r8[1]), .B0(n214), .B1(K_r8[36]), .Y(K10[42])
         );
  AO22X1 U689 ( .A0(n79), .A1(K_r7[15]), .B0(K_r7[22]), .B1(n263), .Y(K9[42])
         );
  AO22X1 U690 ( .A0(n232), .A1(K_r6[15]), .B0(K_r6[22]), .B1(n133), .Y(K8[42])
         );
  AO22X1 U691 ( .A0(n142), .A1(K_r5[36]), .B0(n264), .B1(K_r5[1]), .Y(K7[42])
         );
  AO22X1 U692 ( .A0(n70), .A1(K_r4[50]), .B0(n204), .B1(K_r4[42]), .Y(K6[42])
         );
  AO22X1 U693 ( .A0(n218), .A1(K_r3[28]), .B0(K_r3[9]), .B1(n141), .Y(K5[42])
         );
  AO22X1 U694 ( .A0(n162), .A1(K_r2[14]), .B0(n4), .B1(K_r2[23]), .Y(K4[42])
         );
  AO22X1 U695 ( .A0(n188), .A1(K_r0[45]), .B0(n103), .B1(K_r0[51]), .Y(K2[42])
         );
  AO22X1 U696 ( .A0(n51), .A1(K[31]), .B0(K[38]), .B1(n188), .Y(K1[42]) );
  OAI22X1 U697 ( .A0(n8), .A1(n397), .B0(n165), .B1(n433), .Y(K14[42]) );
  OAI22X1 U698 ( .A0(n160), .A1(n396), .B0(n12), .B1(n432), .Y(K3[42]) );
  AO22X1 U699 ( .A0(K_r14[53]), .A1(n21), .B0(K_r14[46]), .B1(n257), .Y(
        K16[13]) );
  AO22X1 U700 ( .A0(n246), .A1(K_r13[39]), .B0(n34), .B1(K_r13[3]), .Y(K15[13]) );
  AO22X1 U701 ( .A0(n186), .A1(K_r12[25]), .B0(n42), .B1(K_r12[17]), .Y(
        K14[13]) );
  AO22X1 U702 ( .A0(n118), .A1(K_r11[6]), .B0(n272), .B1(K_r11[11]), .Y(
        K13[13]) );
  AO22X1 U703 ( .A0(n185), .A1(K_r10[54]), .B0(n52), .B1(K_r10[20]), .Y(
        K12[13]) );
  AO22X1 U704 ( .A0(n86), .A1(K_r9[34]), .B0(n261), .B1(K_r9[40]), .Y(K11[13])
         );
  AO22X1 U705 ( .A0(n164), .A1(K_r8[26]), .B0(K_r8[48]), .B1(n134), .Y(K10[13]) );
  AO22X1 U706 ( .A0(n195), .A1(K_r7[12]), .B0(K_r7[5]), .B1(n126), .Y(K9[13])
         );
  AO22X1 U707 ( .A0(n132), .A1(K_r6[12]), .B0(K_r6[5]), .B1(n219), .Y(K8[13])
         );
  AO22X1 U708 ( .A0(n75), .A1(K_r5[26]), .B0(K_r5[48]), .B1(n160), .Y(K7[13])
         );
  AO22X1 U709 ( .A0(n254), .A1(K_r4[34]), .B0(n2), .B1(K_r4[40]), .Y(K6[13])
         );
  AO22X1 U710 ( .A0(n66), .A1(K_r3[54]), .B0(n167), .B1(K_r3[20]), .Y(K5[13])
         );
  AO22X1 U711 ( .A0(n169), .A1(K_r2[6]), .B0(n117), .B1(K_r2[11]), .Y(K4[13])
         );
  AO22X1 U712 ( .A0(n65), .A1(K_r1[25]), .B0(n209), .B1(K_r1[17]), .Y(K3[13])
         );
  AO22X1 U713 ( .A0(n55), .A1(K_r0[39]), .B0(n211), .B1(K_r0[3]), .Y(K2[13])
         );
  AO22X1 U714 ( .A0(n264), .A1(K[53]), .B0(K[46]), .B1(n153), .Y(K1[13]) );
  AO22X1 U715 ( .A0(n170), .A1(K_r14[34]), .B0(n117), .B1(K_r14[41]), .Y(
        K16[6]) );
  AO22X1 U716 ( .A0(n37), .A1(K_r13[48]), .B0(n258), .B1(K_r13[27]), .Y(K15[6]) );
  AO22X1 U717 ( .A0(n138), .A1(K_r11[19]), .B0(K_r11[24]), .B1(n196), .Y(
        K13[6]) );
  AO22X1 U718 ( .A0(K_r10[33]), .A1(n22), .B0(K_r10[10]), .B1(n173), .Y(K12[6]) );
  AO22X1 U719 ( .A0(n186), .A1(K_r9[53]), .B0(n25), .B1(K_r9[47]), .Y(K11[6])
         );
  AO22X1 U720 ( .A0(n173), .A1(K_r8[39]), .B0(n104), .B1(K_r8[4]), .Y(K10[6])
         );
  AO22X1 U721 ( .A0(n75), .A1(K_r7[18]), .B0(n205), .B1(K_r7[25]), .Y(K9[6])
         );
  AO22X1 U722 ( .A0(n196), .A1(K_r6[18]), .B0(n134), .B1(K_r6[25]), .Y(K8[6])
         );
  AO22X1 U723 ( .A0(n132), .A1(K_r5[39]), .B0(n233), .B1(K_r5[4]), .Y(K7[6])
         );
  AO22X1 U724 ( .A0(n93), .A1(K_r4[53]), .B0(n245), .B1(K_r4[47]), .Y(K6[6])
         );
  AO22X1 U725 ( .A0(n255), .A1(K_r3[33]), .B0(K_r3[10]), .B1(n143), .Y(K5[6])
         );
  AO22X1 U726 ( .A0(n238), .A1(K_r2[19]), .B0(K_r2[24]), .B1(n125), .Y(K4[6])
         );
  AO22X1 U727 ( .A0(n169), .A1(K_r0[48]), .B0(n107), .B1(K_r0[27]), .Y(K2[6])
         );
  AO22X1 U728 ( .A0(n53), .A1(K[34]), .B0(n212), .B1(K[41]), .Y(K1[6]) );
  OAI22X1 U729 ( .A0(n161), .A1(n425), .B0(n11), .B1(n417), .Y(K14[6]) );
  OAI22X1 U730 ( .A0(n4), .A1(n424), .B0(n165), .B1(n416), .Y(K3[6]) );
  AO22X1 U731 ( .A0(n43), .A1(K_r14[27]), .B0(n269), .B1(K_r14[20]), .Y(K16[7]) );
  AO22X1 U732 ( .A0(n62), .A1(K_r13[34]), .B0(n244), .B1(K_r13[13]), .Y(K15[7]) );
  AO22X1 U733 ( .A0(n137), .A1(K_r11[5]), .B0(n257), .B1(K_r11[10]), .Y(K13[7]) );
  AO22X1 U734 ( .A0(n179), .A1(K_r10[53]), .B0(K_r10[19]), .B1(n138), .Y(
        K12[7]) );
  AO22X1 U735 ( .A0(n186), .A1(K_r9[39]), .B0(K_r9[33]), .B1(n127), .Y(K11[7])
         );
  AO22X1 U736 ( .A0(n84), .A1(K_r8[47]), .B0(n214), .B1(K_r8[25]), .Y(K10[7])
         );
  AO22X1 U737 ( .A0(n75), .A1(K_r7[4]), .B0(n266), .B1(K_r7[11]), .Y(K9[7]) );
  AO22X1 U738 ( .A0(n95), .A1(K_r6[11]), .B0(n213), .B1(K_r6[4]), .Y(K8[7]) );
  AO22X1 U739 ( .A0(n200), .A1(K_r5[47]), .B0(n134), .B1(K_r5[25]), .Y(K7[7])
         );
  AO22X1 U740 ( .A0(K_r4[39]), .A1(n28), .B0(K_r4[33]), .B1(n250), .Y(K6[7])
         );
  AO22X1 U741 ( .A0(K_r3[53]), .A1(n20), .B0(K_r3[19]), .B1(n162), .Y(K5[7])
         );
  AO22X1 U742 ( .A0(n68), .A1(K_r2[10]), .B0(n207), .B1(K_r2[5]), .Y(K4[7]) );
  AO22X1 U743 ( .A0(n174), .A1(K_r0[34]), .B0(n107), .B1(K_r0[13]), .Y(K2[7])
         );
  AO22X1 U744 ( .A0(n179), .A1(K[27]), .B0(n108), .B1(K[20]), .Y(K1[7]) );
  OAI22X1 U745 ( .A0(n160), .A1(n387), .B0(n11), .B1(n407), .Y(K14[7]) );
  OAI22X1 U746 ( .A0(n1), .A1(n386), .B0(n166), .B1(n406), .Y(K3[7]) );
  AO22X1 U747 ( .A0(n47), .A1(K_r14[2]), .B0(K_r14[50]), .B1(n177), .Y(K16[37]) );
  AO22X1 U748 ( .A0(n71), .A1(K_r13[9]), .B0(n208), .B1(K_r13[43]), .Y(K15[37]) );
  AO22X1 U749 ( .A0(n175), .A1(K_r11[15]), .B0(n135), .B1(K_r11[37]), .Y(
        K13[37]) );
  AO22X1 U750 ( .A0(n181), .A1(K_r10[1]), .B0(n47), .B1(K_r10[51]), .Y(K12[37]) );
  AO22X1 U751 ( .A0(n188), .A1(K_r9[42]), .B0(K_r9[38]), .B1(n122), .Y(K11[37]) );
  AO22X1 U752 ( .A0(n80), .A1(K_r8[52]), .B0(n213), .B1(K_r8[28]), .Y(K10[37])
         );
  AO22X1 U753 ( .A0(n192), .A1(K_r7[14]), .B0(K_r7[7]), .B1(n122), .Y(K9[37])
         );
  AO22X1 U754 ( .A0(n98), .A1(K_r6[14]), .B0(K_r6[7]), .B1(n251), .Y(K8[37])
         );
  AO22X1 U755 ( .A0(n202), .A1(K_r5[52]), .B0(n22), .B1(K_r5[28]), .Y(K7[37])
         );
  AO22X1 U756 ( .A0(K_r4[42]), .A1(n19), .B0(K_r4[38]), .B1(n255), .Y(K6[37])
         );
  AO22X1 U757 ( .A0(n57), .A1(K_r3[1]), .B0(n206), .B1(K_r3[51]), .Y(K5[37])
         );
  AO22X1 U758 ( .A0(n72), .A1(K_r2[15]), .B0(n208), .B1(K_r2[37]), .Y(K4[37])
         );
  AO22X1 U759 ( .A0(n186), .A1(K_r0[9]), .B0(n101), .B1(K_r0[43]), .Y(K2[37])
         );
  AO22X1 U760 ( .A0(n176), .A1(K[2]), .B0(K[50]), .B1(n148), .Y(K1[37]) );
  OAI22X1 U761 ( .A0(n9), .A1(n403), .B0(n167), .B1(n409), .Y(K14[37]) );
  OAI22X1 U762 ( .A0(n161), .A1(n402), .B0(n14), .B1(n408), .Y(K3[37]) );
  AO22X1 U763 ( .A0(n55), .A1(K_r14[33]), .B0(n245), .B1(K_r14[26]), .Y(
        K16[15]) );
  AO22X1 U764 ( .A0(K_r13[40]), .A1(n35), .B0(K_r13[19]), .B1(n186), .Y(
        K15[15]) );
  AO22X1 U765 ( .A0(n121), .A1(K_r11[11]), .B0(n266), .B1(K_r11[48]), .Y(
        K13[15]) );
  AO22X1 U766 ( .A0(n98), .A1(K_r10[25]), .B0(K_r10[34]), .B1(n251), .Y(
        K12[15]) );
  AO22X1 U767 ( .A0(n174), .A1(K_r9[20]), .B0(n76), .B1(K_r9[39]), .Y(K11[15])
         );
  AO22X1 U768 ( .A0(n168), .A1(K_r8[6]), .B0(n52), .B1(K_r8[53]), .Y(K10[15])
         );
  AO22X1 U769 ( .A0(n194), .A1(K_r7[17]), .B0(n62), .B1(K_r7[10]), .Y(K9[15])
         );
  AO22X1 U770 ( .A0(n127), .A1(K_r6[17]), .B0(n188), .B1(K_r6[10]), .Y(K8[15])
         );
  AO22X1 U771 ( .A0(n212), .A1(K_r5[53]), .B0(n143), .B1(K_r5[6]), .Y(K7[15])
         );
  AO22X1 U772 ( .A0(n47), .A1(K_r4[20]), .B0(n205), .B1(K_r4[39]), .Y(K6[15])
         );
  AO22X1 U773 ( .A0(n228), .A1(K_r3[25]), .B0(K_r3[34]), .B1(n127), .Y(K5[15])
         );
  AO22X1 U774 ( .A0(n171), .A1(K_r2[11]), .B0(n116), .B1(K_r2[48]), .Y(K4[15])
         );
  AO22X1 U775 ( .A0(n180), .A1(K_r0[40]), .B0(K_r0[19]), .B1(n140), .Y(K2[15])
         );
  AO22X1 U776 ( .A0(n215), .A1(K[33]), .B0(n118), .B1(K[26]), .Y(K1[15]) );
  OAI22X1 U777 ( .A0(n4), .A1(n425), .B0(n162), .B1(n379), .Y(K14[15]) );
  OAI22X1 U778 ( .A0(n158), .A1(n424), .B0(n9), .B1(n378), .Y(K3[15]) );
  AO22X1 U779 ( .A0(n39), .A1(K_r14[16]), .B0(n212), .B1(K_r14[9]), .Y(K16[43]) );
  AO22X1 U780 ( .A0(n60), .A1(K_r13[23]), .B0(K_r13[2]), .B1(n161), .Y(K15[43]) );
  AO22X1 U781 ( .A0(K_r11[51]), .A1(n25), .B0(K_r11[29]), .B1(n203), .Y(
        K13[43]) );
  AO22X1 U782 ( .A0(n180), .A1(K_r10[15]), .B0(n29), .B1(K_r10[38]), .Y(
        K12[43]) );
  AO22X1 U783 ( .A0(n94), .A1(K_r9[52]), .B0(n232), .B1(K_r9[1]), .Y(K11[43])
         );
  AO22X1 U784 ( .A0(n82), .A1(K_r8[7]), .B0(n214), .B1(K_r8[42]), .Y(K10[43])
         );
  AO22X1 U785 ( .A0(n191), .A1(K_r7[28]), .B0(n95), .B1(K_r7[21]), .Y(K9[43])
         );
  AO22X1 U786 ( .A0(n97), .A1(K_r6[28]), .B0(n208), .B1(K_r6[21]), .Y(K8[43])
         );
  AO22X1 U787 ( .A0(n201), .A1(K_r5[7]), .B0(n97), .B1(K_r5[42]), .Y(K7[43])
         );
  AO22X1 U788 ( .A0(n85), .A1(K_r4[1]), .B0(n243), .B1(K_r4[52]), .Y(K6[43])
         );
  AO22X1 U789 ( .A0(n53), .A1(K_r3[15]), .B0(n206), .B1(K_r3[38]), .Y(K5[43])
         );
  AO22X1 U790 ( .A0(n164), .A1(K_r2[51]), .B0(K_r2[29]), .B1(n124), .Y(K4[43])
         );
  AO22X1 U791 ( .A0(n188), .A1(K_r0[23]), .B0(K_r0[2]), .B1(n129), .Y(K2[43])
         );
  AO22X1 U792 ( .A0(n177), .A1(K[16]), .B0(n109), .B1(K[9]), .Y(K1[43]) );
  OAI22X1 U793 ( .A0(n2), .A1(n393), .B0(n166), .B1(n397), .Y(K14[43]) );
  OAI22X1 U794 ( .A0(n162), .A1(n392), .B0(n9), .B1(n396), .Y(K3[43]) );
  AO22X1 U795 ( .A0(n203), .A1(K_r14[21]), .B0(n119), .B1(K_r14[28]), .Y(
        K16[48]) );
  AO22X1 U796 ( .A0(n197), .A1(K_r13[14]), .B0(K_r13[35]), .B1(n152), .Y(
        K15[48]) );
  AO22X1 U797 ( .A0(n180), .A1(K_r11[45]), .B0(K_r11[8]), .B1(n143), .Y(
        K13[48]) );
  AO22X1 U798 ( .A0(n76), .A1(K_r10[22]), .B0(n271), .B1(K_r10[31]), .Y(
        K12[48]) );
  AO22X1 U799 ( .A0(n186), .A1(K_r9[44]), .B0(n136), .B1(K_r9[36]), .Y(K11[48]) );
  AO22X1 U800 ( .A0(n172), .A1(K_r8[30]), .B0(n66), .B1(K_r8[50]), .Y(K10[48])
         );
  AO22X1 U801 ( .A0(n77), .A1(K_r7[9]), .B0(n241), .B1(K_r7[16]), .Y(K9[48])
         );
  AO22X1 U802 ( .A0(n196), .A1(K_r6[9]), .B0(n56), .B1(K_r6[16]), .Y(K8[48])
         );
  AO22X1 U803 ( .A0(n133), .A1(K_r5[30]), .B0(n261), .B1(K_r5[50]), .Y(K7[48])
         );
  AO22X1 U804 ( .A0(n37), .A1(K_r4[44]), .B0(n259), .B1(K_r4[36]), .Y(K6[48])
         );
  AO22X1 U805 ( .A0(n242), .A1(K_r3[22]), .B0(n10), .B1(K_r3[31]), .Y(K5[48])
         );
  AO22X1 U806 ( .A0(n69), .A1(K_r2[45]), .B0(K_r2[8]), .B1(n247), .Y(K4[48])
         );
  AO22X1 U807 ( .A0(n63), .A1(K_r0[14]), .B0(K_r0[35]), .B1(n161), .Y(K2[48])
         );
  AO22X1 U808 ( .A0(n53), .A1(K[21]), .B0(n212), .B1(K[28]), .Y(K1[48]) );
  OAI22X1 U809 ( .A0(n162), .A1(n385), .B0(n16), .B1(n433), .Y(K14[48]) );
  OAI22X1 U810 ( .A0(n4), .A1(n384), .B0(n166), .B1(n432), .Y(K3[48]) );
  AO22X1 U811 ( .A0(n84), .A1(K_r14[20]), .B0(n244), .B1(K_r14[13]), .Y(
        K16[24]) );
  AO22X1 U812 ( .A0(n32), .A1(K_r13[27]), .B0(n213), .B1(K_r13[6]), .Y(K15[24]) );
  AO22X1 U813 ( .A0(n172), .A1(K_r12[17]), .B0(K_r12[41]), .B1(n144), .Y(
        K14[24]) );
  AO22X1 U814 ( .A0(n123), .A1(K_r11[55]), .B0(n265), .B1(K_r11[3]), .Y(
        K13[24]) );
  AO22X1 U815 ( .A0(n100), .A1(K_r10[12]), .B0(n251), .B1(K_r10[46]), .Y(
        K12[24]) );
  AO22X1 U816 ( .A0(n189), .A1(K_r9[32]), .B0(n60), .B1(K_r9[26]), .Y(K11[24])
         );
  AO22X1 U817 ( .A0(n168), .A1(K_r8[18]), .B0(K_r8[40]), .B1(n130), .Y(K10[24]) );
  AO22X1 U818 ( .A0(n193), .A1(K_r7[4]), .B0(n74), .B1(K_r7[54]), .Y(K9[24])
         );
  AO22X1 U819 ( .A0(n64), .A1(K_r6[4]), .B0(n199), .B1(K_r6[54]), .Y(K8[24])
         );
  AO22X1 U820 ( .A0(n124), .A1(K_r5[18]), .B0(K_r5[40]), .B1(n249), .Y(K7[24])
         );
  AO22X1 U821 ( .A0(n45), .A1(K_r4[32]), .B0(n205), .B1(K_r4[26]), .Y(K6[24])
         );
  AO22X1 U822 ( .A0(n217), .A1(K_r3[12]), .B0(n154), .B1(K_r3[46]), .Y(K5[24])
         );
  AO22X1 U823 ( .A0(n172), .A1(K_r2[55]), .B0(n118), .B1(K_r2[3]), .Y(K4[24])
         );
  AO22X1 U824 ( .A0(n66), .A1(K_r1[17]), .B0(K_r1[41]), .B1(n252), .Y(K3[24])
         );
  AO22X1 U825 ( .A0(n183), .A1(K_r0[27]), .B0(n104), .B1(K_r0[6]), .Y(K2[24])
         );
  AO22X1 U826 ( .A0(n181), .A1(K[20]), .B0(n113), .B1(K[13]), .Y(K1[24]) );
  AO22X1 U827 ( .A0(K_r14[19]), .A1(n25), .B0(K_r14[12]), .B1(n243), .Y(
        K16[12]) );
  AO22X1 U828 ( .A0(n223), .A1(K_r13[5]), .B0(n31), .B1(K_r13[26]), .Y(K15[12]) );
  AO22X1 U829 ( .A0(n126), .A1(K_r11[54]), .B0(n269), .B1(K_r11[34]), .Y(
        K13[12]) );
  AO22X1 U830 ( .A0(n185), .A1(K_r10[20]), .B0(K_r10[11]), .B1(n132), .Y(
        K12[12]) );
  AO22X1 U831 ( .A0(n85), .A1(K_r9[25]), .B0(n262), .B1(K_r9[6]), .Y(K11[12])
         );
  AO22X1 U832 ( .A0(n75), .A1(K_r8[39]), .B0(n211), .B1(K_r8[17]), .Y(K10[12])
         );
  AO22X1 U833 ( .A0(n195), .A1(K_r7[3]), .B0(K_r7[53]), .B1(n126), .Y(K9[12])
         );
  AO22X1 U834 ( .A0(n130), .A1(K_r6[3]), .B0(K_r6[53]), .B1(n164), .Y(K8[12])
         );
  AO22X1 U835 ( .A0(n239), .A1(K_r5[39]), .B0(n110), .B1(K_r5[17]), .Y(K7[12])
         );
  AO22X1 U836 ( .A0(n157), .A1(K_r4[25]), .B0(n144), .B1(K_r4[6]), .Y(K6[12])
         );
  AO22X1 U837 ( .A0(K_r3[20]), .A1(n32), .B0(K_r3[11]), .B1(n242), .Y(K5[12])
         );
  AO22X1 U838 ( .A0(n170), .A1(K_r2[54]), .B0(n114), .B1(K_r2[34]), .Y(K4[12])
         );
  AO22X1 U839 ( .A0(n55), .A1(K_r0[5]), .B0(n212), .B1(K_r0[26]), .Y(K2[12])
         );
  AO22X1 U840 ( .A0(n194), .A1(K[19]), .B0(K[12]), .B1(n154), .Y(K1[12]) );
  OAI22X1 U841 ( .A0(n1), .A1(n387), .B0(n163), .B1(n395), .Y(K14[12]) );
  OAI22X1 U842 ( .A0(n157), .A1(n386), .B0(n16), .B1(n394), .Y(K3[12]) );
  AO22X1 U843 ( .A0(n192), .A1(K_r14[55]), .B0(K_r14[5]), .B1(n154), .Y(
        K16[18]) );
  AO22X1 U844 ( .A0(n125), .A1(K_r13[12]), .B0(n214), .B1(K_r13[48]), .Y(
        K15[18]) );
  AO22X1 U845 ( .A0(n188), .A1(K_r12[34]), .B0(n41), .B1(K_r12[26]), .Y(
        K14[18]) );
  AO22X1 U846 ( .A0(K_r11[40]), .A1(n22), .B0(K_r11[20]), .B1(n172), .Y(
        K13[18]) );
  AO22X1 U847 ( .A0(n184), .A1(K_r10[6]), .B0(n101), .B1(K_r10[54]), .Y(
        K12[18]) );
  AO22X1 U848 ( .A0(n174), .A1(K_r9[17]), .B0(n78), .B1(K_r9[11]), .Y(K11[18])
         );
  AO22X1 U849 ( .A0(n76), .A1(K_r8[25]), .B0(n240), .B1(K_r8[3]), .Y(K10[18])
         );
  AO22X1 U850 ( .A0(n91), .A1(K_r7[39]), .B0(K_r7[46]), .B1(n240), .Y(K9[18])
         );
  AO22X1 U851 ( .A0(n199), .A1(K_r6[39]), .B0(K_r6[46]), .B1(n139), .Y(K8[18])
         );
  AO22X1 U852 ( .A0(n214), .A1(K_r5[25]), .B0(n147), .B1(K_r5[3]), .Y(K7[18])
         );
  AO22X1 U853 ( .A0(n47), .A1(K_r4[17]), .B0(n205), .B1(K_r4[11]), .Y(K6[18])
         );
  AO22X1 U854 ( .A0(n64), .A1(K_r3[6]), .B0(n165), .B1(K_r3[54]), .Y(K5[18])
         );
  AO22X1 U855 ( .A0(n171), .A1(K_r2[40]), .B0(K_r2[20]), .B1(n125), .Y(K4[18])
         );
  AO22X1 U856 ( .A0(n239), .A1(K_r1[26]), .B0(n109), .B1(K_r1[34]), .Y(K3[18])
         );
  AO22X1 U857 ( .A0(n180), .A1(K_r0[12]), .B0(n106), .B1(K_r0[48]), .Y(K2[18])
         );
  AO22X1 U858 ( .A0(n46), .A1(K[55]), .B0(K[5]), .B1(n194), .Y(K1[18]) );
  OAI22X1 U859 ( .A0(n159), .A1(n383), .B0(n18), .B1(n431), .Y(K14[36]) );
  OAI22X1 U860 ( .A0(n6), .A1(n382), .B0(n164), .B1(n430), .Y(K3[36]) );
  AO22X1 U861 ( .A0(n51), .A1(K_r14[30]), .B0(n263), .B1(K_r14[23]), .Y(
        K16[36]) );
  AO22X1 U862 ( .A0(n200), .A1(K_r13[16]), .B0(n37), .B1(K_r13[37]), .Y(
        K15[36]) );
  AO22X1 U863 ( .A0(n142), .A1(K_r11[38]), .B0(n271), .B1(K_r11[43]), .Y(
        K13[36]) );
  AO22X1 U864 ( .A0(n181), .A1(K_r10[29]), .B0(K_r10[52]), .B1(n136), .Y(
        K12[36]) );
  AO22X1 U865 ( .A0(n92), .A1(K_r9[7]), .B0(n248), .B1(K_r9[15]), .Y(K11[36])
         );
  AO22X1 U866 ( .A0(n171), .A1(K_r8[1]), .B0(K_r8[21]), .B1(n128), .Y(K10[36])
         );
  AO22X1 U867 ( .A0(n192), .A1(K_r7[42]), .B0(n38), .B1(K_r7[35]), .Y(K9[36])
         );
  AO22X1 U868 ( .A0(n99), .A1(K_r6[42]), .B0(n162), .B1(K_r6[35]), .Y(K8[36])
         );
  AO22X1 U869 ( .A0(n29), .A1(K_r5[1]), .B0(K_r5[21]), .B1(n168), .Y(K7[36])
         );
  AO22X1 U870 ( .A0(n180), .A1(K_r4[7]), .B0(n152), .B1(K_r4[15]), .Y(K6[36])
         );
  AO22X1 U871 ( .A0(n58), .A1(K_r3[29]), .B0(K_r3[52]), .B1(n248), .Y(K5[36])
         );
  AO22X1 U872 ( .A0(n231), .A1(K_r2[38]), .B0(n45), .B1(K_r2[43]), .Y(K4[36])
         );
  AO22X1 U873 ( .A0(n61), .A1(K_r0[16]), .B0(n210), .B1(K_r0[37]), .Y(K2[36])
         );
  AO22X1 U874 ( .A0(n175), .A1(K[30]), .B0(n111), .B1(K[23]), .Y(K1[36]) );
  CLKINVX1 U875 ( .A(K_r12[51]), .Y(n383) );
  CLKINVX1 U876 ( .A(K_r1[51]), .Y(n382) );
  CLKINVX1 U877 ( .A(K_r12[49]), .Y(n385) );
  CLKINVX1 U878 ( .A(K_r12[45]), .Y(n391) );
  CLKINVX1 U879 ( .A(K_r12[5]), .Y(n425) );
  CLKINVX1 U880 ( .A(K_r12[48]), .Y(n387) );
  CLKINVX1 U881 ( .A(K_r1[49]), .Y(n384) );
  CLKINVX1 U882 ( .A(K_r1[45]), .Y(n390) );
  CLKINVX1 U883 ( .A(K_r1[5]), .Y(n424) );
  CLKINVX1 U884 ( .A(K_r1[48]), .Y(n386) );
  CLKINVX1 U885 ( .A(K_r12[3]), .Y(n429) );
  CLKINVX1 U886 ( .A(K_r1[3]), .Y(n428) );
  CLKINVX1 U887 ( .A(K_r12[53]), .Y(n381) );
  CLKINVX1 U888 ( .A(K_r12[8]), .Y(n423) );
  CLKINVX1 U889 ( .A(K_r1[53]), .Y(n380) );
  CLKINVX1 U890 ( .A(K_r1[8]), .Y(n422) );
  CLKINVX1 U891 ( .A(K_r12[37]), .Y(n397) );
  CLKINVX1 U892 ( .A(K_r12[43]), .Y(n393) );
  CLKINVX1 U893 ( .A(K_r12[32]), .Y(n401) );
  CLKINVX1 U894 ( .A(K_r12[29]), .Y(n403) );
  CLKINVX1 U895 ( .A(K_r12[54]), .Y(n379) );
  CLKINVX1 U896 ( .A(K_r12[40]), .Y(n395) );
  CLKINVX1 U897 ( .A(K_r1[37]), .Y(n396) );
  CLKINVX1 U898 ( .A(K_r1[43]), .Y(n392) );
  CLKINVX1 U899 ( .A(K_r1[32]), .Y(n400) );
  CLKINVX1 U900 ( .A(K_r1[29]), .Y(n402) );
  CLKINVX1 U901 ( .A(K_r1[54]), .Y(n378) );
  CLKINVX1 U902 ( .A(K_r1[40]), .Y(n394) );
  CLKINVX1 U903 ( .A(K_r12[46]), .Y(n389) );
  CLKINVX1 U904 ( .A(K_r12[20]), .Y(n411) );
  CLKINVX1 U905 ( .A(K_r1[46]), .Y(n388) );
  CLKINVX1 U906 ( .A(K_r1[20]), .Y(n410) );
  CLKINVX1 U907 ( .A(K_r12[4]), .Y(n427) );
  CLKINVX1 U908 ( .A(K_r12[19]), .Y(n413) );
  CLKINVX1 U909 ( .A(K_r12[35]), .Y(n399) );
  CLKINVX1 U910 ( .A(K_r12[27]), .Y(n405) );
  CLKINVX1 U911 ( .A(K_r1[4]), .Y(n426) );
  CLKINVX1 U912 ( .A(K_r1[19]), .Y(n412) );
  CLKINVX1 U913 ( .A(K_r1[35]), .Y(n398) );
  CLKINVX1 U914 ( .A(K_r1[27]), .Y(n404) );
  CLKINVX1 U915 ( .A(K_r12[2]), .Y(n431) );
  CLKINVX1 U916 ( .A(K_r1[2]), .Y(n430) );
  CLKINVX1 U917 ( .A(K_r12[0]), .Y(n433) );
  CLKINVX1 U918 ( .A(K_r12[24]), .Y(n407) );
  CLKINVX1 U919 ( .A(K_r12[14]), .Y(n415) );
  CLKINVX1 U920 ( .A(K_r12[23]), .Y(n409) );
  CLKINVX1 U921 ( .A(K_r1[0]), .Y(n432) );
  CLKINVX1 U922 ( .A(K_r1[24]), .Y(n406) );
  CLKINVX1 U923 ( .A(K_r1[14]), .Y(n414) );
  CLKINVX1 U924 ( .A(K_r1[23]), .Y(n408) );
  CLKINVX1 U925 ( .A(K_r12[12]), .Y(n419) );
  CLKINVX1 U926 ( .A(K_r1[12]), .Y(n418) );
  CLKINVX1 U927 ( .A(K_r12[11]), .Y(n421) );
  CLKINVX1 U928 ( .A(K_r1[11]), .Y(n420) );
  CLKINVX1 U929 ( .A(K_r12[13]), .Y(n417) );
  CLKINVX1 U930 ( .A(K_r1[13]), .Y(n416) );
  AO22X1 U931 ( .A0(n195), .A1(K_r14[4]), .B0(K_r14[11]), .B1(n156), .Y(K16[2]) );
  AO22X1 U932 ( .A0(n40), .A1(K_r13[18]), .B0(n159), .B1(K_r13[54]), .Y(K15[2]) );
  OAI22X1 U933 ( .A0(n2), .A1(n395), .B0(n168), .B1(n401), .Y(K14[2]) );
  AO22X1 U934 ( .A0(n176), .A1(K_r11[26]), .B0(n81), .B1(K_r11[46]), .Y(K13[2]) );
  AO22X1 U935 ( .A0(n39), .A1(K_r10[3]), .B0(n266), .B1(K_r10[12]), .Y(K12[2])
         );
  AO22X1 U936 ( .A0(n189), .A1(K_r9[55]), .B0(n7), .B1(K_r9[17]), .Y(K11[2])
         );
  AO22X1 U937 ( .A0(K_r8[6]), .A1(n31), .B0(K_r8[41]), .B1(n157), .Y(K10[2])
         );
  AO22X1 U938 ( .A0(n84), .A1(K_r7[20]), .B0(K_r7[27]), .B1(n246), .Y(K9[2])
         );
  AO22X1 U939 ( .A0(n198), .A1(K_r6[20]), .B0(K_r6[27]), .B1(n136), .Y(K8[2])
         );
  AO22X1 U940 ( .A0(n203), .A1(K_r5[6]), .B0(K_r5[41]), .B1(n147), .Y(K7[2])
         );
  AO22X1 U941 ( .A0(n40), .A1(K_r4[55]), .B0(n204), .B1(K_r4[17]), .Y(K6[2])
         );
  AO22X1 U942 ( .A0(n189), .A1(K_r3[3]), .B0(n144), .B1(K_r3[12]), .Y(K5[2])
         );
  AO22X1 U943 ( .A0(n41), .A1(K_r2[26]), .B0(n208), .B1(K_r2[46]), .Y(K4[2])
         );
  OAI22X1 U944 ( .A0(n160), .A1(n394), .B0(n12), .B1(n400), .Y(K3[2]) );
  AO22X1 U945 ( .A0(n184), .A1(K_r0[18]), .B0(n103), .B1(K_r0[54]), .Y(K2[2])
         );
  AO22X1 U946 ( .A0(K[4]), .A1(n20), .B0(K[11]), .B1(n176), .Y(K1[2]) );
  AO22X1 U947 ( .A0(n68), .A1(K_r14[9]), .B0(n162), .B1(K_r14[2]), .Y(K16[34])
         );
  AO22X1 U948 ( .A0(n201), .A1(K_r13[50]), .B0(n96), .B1(K_r13[16]), .Y(
        K15[34]) );
  AO22X1 U949 ( .A0(n119), .A1(K_r12[30]), .B0(K_r12[36]), .B1(n159), .Y(
        K14[34]) );
  AO22X1 U950 ( .A0(n130), .A1(K_r11[44]), .B0(n269), .B1(K_r11[22]), .Y(
        K13[34]) );
  AO22X1 U951 ( .A0(n21), .A1(K_r10[31]), .B0(n249), .B1(K_r10[8]), .Y(K12[34]) );
  AO22X1 U952 ( .A0(n91), .A1(K_r9[45]), .B0(K_r9[49]), .B1(n213), .Y(K11[34])
         );
  AO22X1 U953 ( .A0(n170), .A1(K_r8[35]), .B0(n80), .B1(K_r8[0]), .Y(K10[34])
         );
  AO22X1 U954 ( .A0(n192), .A1(K_r7[21]), .B0(decrypt), .B1(K_r7[14]), .Y(
        K9[34]) );
  AO22X1 U955 ( .A0(n37), .A1(K_r6[21]), .B0(n205), .B1(K_r6[14]), .Y(K8[34])
         );
  AO22X1 U956 ( .A0(n101), .A1(K_r5[35]), .B0(n234), .B1(K_r5[0]), .Y(K7[34])
         );
  AO22X1 U957 ( .A0(n182), .A1(K_r4[45]), .B0(K_r4[49]), .B1(n134), .Y(K6[34])
         );
  AO22X1 U958 ( .A0(n190), .A1(K_r3[31]), .B0(n102), .B1(K_r3[8]), .Y(K5[34])
         );
  AO22X1 U959 ( .A0(n221), .A1(K_r2[44]), .B0(n149), .B1(K_r2[22]), .Y(K4[34])
         );
  AO22X1 U960 ( .A0(n166), .A1(K_r1[30]), .B0(K_r1[36]), .B1(n121), .Y(K3[34])
         );
  AO22X1 U961 ( .A0(n60), .A1(K_r0[50]), .B0(n210), .B1(K_r0[16]), .Y(K2[34])
         );
  AO22X1 U962 ( .A0(n175), .A1(K[9]), .B0(n112), .B1(K[2]), .Y(K1[34]) );
  AO22X1 U963 ( .A0(K_r14[25]), .A1(n21), .B0(K_r14[18]), .B1(n187), .Y(
        K16[14]) );
  AO22X1 U964 ( .A0(n183), .A1(K_r13[11]), .B0(K_r13[32]), .B1(n135), .Y(
        K15[14]) );
  OAI22X1 U965 ( .A0(n3), .A1(n379), .B0(n164), .B1(n389), .Y(K14[14]) );
  AO22X1 U966 ( .A0(n150), .A1(K_r11[3]), .B0(n260), .B1(K_r11[40]), .Y(
        K13[14]) );
  AO22X1 U967 ( .A0(n185), .A1(K_r10[26]), .B0(n82), .B1(K_r10[17]), .Y(
        K12[14]) );
  AO22X1 U968 ( .A0(n86), .A1(K_r9[6]), .B0(n240), .B1(K_r9[12]), .Y(K11[14])
         );
  AO22X1 U969 ( .A0(n169), .A1(K_r8[55]), .B0(n90), .B1(K_r8[20]), .Y(K10[14])
         );
  AO22X1 U970 ( .A0(n195), .A1(K_r7[41]), .B0(K_r7[34]), .B1(n126), .Y(K9[14])
         );
  AO22X1 U971 ( .A0(K_r6[41]), .A1(n18), .B0(K_r6[34]), .B1(n267), .Y(K8[14])
         );
  AO22X1 U972 ( .A0(n83), .A1(K_r5[55]), .B0(n238), .B1(K_r5[20]), .Y(K7[14])
         );
  AO22X1 U973 ( .A0(n192), .A1(K_r4[6]), .B0(n147), .B1(K_r4[12]), .Y(K6[14])
         );
  AO22X1 U974 ( .A0(n66), .A1(K_r3[26]), .B0(n238), .B1(K_r3[17]), .Y(K5[14])
         );
  AO22X1 U975 ( .A0(n228), .A1(K_r2[3]), .B0(n115), .B1(K_r2[40]), .Y(K4[14])
         );
  OAI22X1 U976 ( .A0(n157), .A1(n378), .B0(n15), .B1(n388), .Y(K3[14]) );
  AO22X1 U977 ( .A0(n56), .A1(K_r0[11]), .B0(K_r0[32]), .B1(n236), .Y(K2[14])
         );
  AO22X1 U978 ( .A0(n217), .A1(K[25]), .B0(K[18]), .B1(n151), .Y(K1[14]) );
  AO22X1 U979 ( .A0(n201), .A1(K_r14[37]), .B0(n117), .B1(K_r14[44]), .Y(
        K16[45]) );
  AO22X1 U980 ( .A0(n63), .A1(K_r13[51]), .B0(n230), .B1(K_r13[30]), .Y(
        K15[45]) );
  AO22X1 U981 ( .A0(K_r12[38]), .A1(n31), .B0(K_r12[16]), .B1(n192), .Y(
        K14[45]) );
  AO22X1 U982 ( .A0(n178), .A1(K_r11[2]), .B0(n72), .B1(K_r11[52]), .Y(K13[45]) );
  AO22X1 U983 ( .A0(K_r10[7]), .A1(n23), .B0(K_r10[43]), .B1(n247), .Y(K12[45]) );
  AO22X1 U984 ( .A0(n187), .A1(K_r9[29]), .B0(n137), .B1(K_r9[21]), .Y(K11[45]) );
  AO22X1 U985 ( .A0(n172), .A1(K_r8[15]), .B0(n87), .B1(K_r8[35]), .Y(K10[45])
         );
  AO22X1 U986 ( .A0(n78), .A1(K_r7[49]), .B0(n245), .B1(K_r7[1]), .Y(K9[45])
         );
  AO22X1 U987 ( .A0(n196), .A1(K_r6[49]), .B0(n101), .B1(K_r6[1]), .Y(K8[45])
         );
  AO22X1 U988 ( .A0(n106), .A1(K_r5[15]), .B0(n267), .B1(K_r5[35]), .Y(K7[45])
         );
  AO22X1 U989 ( .A0(n54), .A1(K_r4[29]), .B0(n258), .B1(K_r4[21]), .Y(K6[45])
         );
  AO22X1 U990 ( .A0(n216), .A1(K_r3[7]), .B0(K_r3[43]), .B1(n142), .Y(K5[45])
         );
  AO22X1 U991 ( .A0(n70), .A1(K_r2[2]), .B0(n207), .B1(K_r2[52]), .Y(K4[45])
         );
  AO22X1 U992 ( .A0(n165), .A1(K_r1[38]), .B0(K_r1[16]), .B1(n122), .Y(K3[45])
         );
  AO22X1 U993 ( .A0(n188), .A1(K_r0[51]), .B0(n105), .B1(K_r0[30]), .Y(K2[45])
         );
  AO22X1 U994 ( .A0(n52), .A1(K[37]), .B0(n212), .B1(K[44]), .Y(K1[45]) );
  AO22X1 U995 ( .A0(n39), .A1(K_r14[29]), .B0(n262), .B1(K_r14[22]), .Y(
        K16[32]) );
  AO22X1 U996 ( .A0(n201), .A1(K_r13[15]), .B0(K_r13[36]), .B1(n149), .Y(
        K15[32]) );
  AO22X1 U997 ( .A0(n33), .A1(K_r12[50]), .B0(n241), .B1(K_r12[1]), .Y(K14[32]) );
  AO22X1 U998 ( .A0(n139), .A1(K_r11[9]), .B0(n266), .B1(K_r11[42]), .Y(
        K13[32]) );
  AO22X1 U999 ( .A0(n43), .A1(K_r10[23]), .B0(n221), .B1(K_r10[28]), .Y(
        K12[32]) );
  AO22X1 U1000 ( .A0(n90), .A1(K_r9[37]), .B0(n250), .B1(K_r9[14]), .Y(K11[32]) );
  AO22X1 U1001 ( .A0(n170), .A1(K_r8[0]), .B0(K_r8[51]), .B1(n129), .Y(K10[32]) );
  AO22X1 U1002 ( .A0(n192), .A1(K_r7[45]), .B0(n56), .B1(K_r7[38]), .Y(K9[32])
         );
  AO22X1 U1003 ( .A0(n40), .A1(K_r6[45]), .B0(n204), .B1(K_r6[38]), .Y(K8[32])
         );
  AO22X1 U1004 ( .A0(n109), .A1(K_r5[0]), .B0(K_r5[51]), .B1(n157), .Y(K7[32])
         );
  AO22X1 U1005 ( .A0(n261), .A1(K_r4[37]), .B0(n153), .B1(K_r4[14]), .Y(K6[32]) );
  AO22X1 U1006 ( .A0(n191), .A1(K_r3[23]), .B0(n18), .B1(K_r3[28]), .Y(K5[32])
         );
  AO22X1 U1007 ( .A0(n174), .A1(K_r2[9]), .B0(n111), .B1(K_r2[42]), .Y(K4[32])
         );
  AO22X1 U1008 ( .A0(n168), .A1(K_r1[50]), .B0(n110), .B1(K_r1[1]), .Y(K3[32])
         );
  AO22X1 U1009 ( .A0(n60), .A1(K_r0[15]), .B0(K_r0[36]), .B1(n244), .Y(K2[32])
         );
  AO22X1 U1010 ( .A0(n175), .A1(K[29]), .B0(n112), .B1(K[22]), .Y(K1[32]) );
  AO22X1 U1011 ( .A0(n198), .A1(K_r14[30]), .B0(n101), .B1(K_r14[37]), .Y(
        K16[38]) );
  AO22X1 U1012 ( .A0(n37), .A1(K_r13[44]), .B0(n243), .B1(K_r13[23]), .Y(
        K15[38]) );
  AO22X1 U1013 ( .A0(n227), .A1(K_r12[9]), .B0(n30), .B1(K_r12[31]), .Y(
        K14[38]) );
  AO22X1 U1014 ( .A0(n139), .A1(K_r11[45]), .B0(K_r11[50]), .B1(n195), .Y(
        K13[38]) );
  AO22X1 U1015 ( .A0(n181), .A1(K_r10[36]), .B0(n65), .B1(K_r10[0]), .Y(
        K12[38]) );
  AO22X1 U1016 ( .A0(n92), .A1(K_r9[14]), .B0(n249), .B1(K_r9[22]), .Y(K11[38]) );
  AO22X1 U1017 ( .A0(n80), .A1(K_r8[28]), .B0(K_r8[8]), .B1(n238), .Y(K10[38])
         );
  AO22X1 U1018 ( .A0(n81), .A1(K_r7[42]), .B0(n243), .B1(K_r7[49]), .Y(K9[38])
         );
  AO22X1 U1019 ( .A0(n197), .A1(K_r6[42]), .B0(n15), .B1(K_r6[49]), .Y(K8[38])
         );
  AO22X1 U1020 ( .A0(n202), .A1(K_r5[28]), .B0(K_r5[8]), .B1(n144), .Y(K7[38])
         );
  AO22X1 U1021 ( .A0(n172), .A1(K_r4[14]), .B0(n69), .B1(K_r4[22]), .Y(K6[38])
         );
  AO22X1 U1022 ( .A0(n57), .A1(K_r3[36]), .B0(n206), .B1(K_r3[0]), .Y(K5[38])
         );
  AO22X1 U1023 ( .A0(n163), .A1(K_r2[45]), .B0(K_r2[50]), .B1(n131), .Y(K4[38]) );
  AO22X1 U1024 ( .A0(n168), .A1(K_r1[31]), .B0(n111), .B1(K_r1[9]), .Y(K3[38])
         );
  AO22X1 U1025 ( .A0(n187), .A1(K_r0[44]), .B0(n113), .B1(K_r0[23]), .Y(K2[38]) );
  AO22X1 U1026 ( .A0(n50), .A1(K[30]), .B0(n212), .B1(K[37]), .Y(K1[38]) );
  AO22X1 U1027 ( .A0(n39), .A1(K_r14[0]), .B0(n248), .B1(K_r14[52]), .Y(
        K16[40]) );
  AO22X1 U1028 ( .A0(n53), .A1(K_r13[7]), .B0(n227), .B1(K_r13[45]), .Y(
        K15[40]) );
  AO22X1 U1029 ( .A0(n229), .A1(K_r12[31]), .B0(K_r12[21]), .B1(n146), .Y(
        K14[40]) );
  AO22X1 U1030 ( .A0(n190), .A1(K_r11[44]), .B0(n81), .B1(K_r11[35]), .Y(
        K13[40]) );
  AO22X1 U1031 ( .A0(n181), .A1(K_r10[30]), .B0(K_r10[49]), .B1(n137), .Y(
        K12[40]) );
  AO22X1 U1032 ( .A0(n187), .A1(K_r9[16]), .B0(n120), .B1(K_r9[8]), .Y(K11[40]) );
  AO22X1 U1033 ( .A0(n81), .A1(K_r8[22]), .B0(n214), .B1(K_r8[2]), .Y(K10[40])
         );
  AO22X1 U1034 ( .A0(n191), .A1(K_r7[43]), .B0(n91), .B1(K_r7[36]), .Y(K9[40])
         );
  AO22X1 U1035 ( .A0(n97), .A1(K_r6[43]), .B0(n206), .B1(K_r6[36]), .Y(K8[40])
         );
  AO22X1 U1036 ( .A0(n202), .A1(K_r5[22]), .B0(n58), .B1(K_r5[2]), .Y(K7[40])
         );
  AO22X1 U1037 ( .A0(n73), .A1(K_r4[16]), .B0(n204), .B1(K_r4[8]), .Y(K6[40])
         );
  AO22X1 U1038 ( .A0(n54), .A1(K_r3[30]), .B0(K_r3[49]), .B1(n250), .Y(K5[40])
         );
  AO22X1 U1039 ( .A0(n71), .A1(K_r2[44]), .B0(n207), .B1(K_r2[35]), .Y(K4[40])
         );
  AO22X1 U1040 ( .A0(K_r1[31]), .A1(n34), .B0(K_r1[21]), .B1(n251), .Y(K3[40])
         );
  AO22X1 U1041 ( .A0(n62), .A1(K_r0[45]), .B0(n210), .B1(K_r0[7]), .Y(K2[40])
         );
  AO22X1 U1042 ( .A0(n177), .A1(K[0]), .B0(n109), .B1(K[52]), .Y(K1[40]) );
  AO22X1 U1043 ( .A0(n184), .A1(K_r14[53]), .B0(K_r14[3]), .B1(n154), .Y(
        K16[4]) );
  AO22X1 U1044 ( .A0(n59), .A1(K_r13[10]), .B0(n263), .B1(K_r13[46]), .Y(
        K15[4]) );
  OAI22X1 U1045 ( .A0(decrypt), .A1(n401), .B0(n164), .B1(n407), .Y(K14[4]) );
  AO22X1 U1046 ( .A0(n180), .A1(K_r11[18]), .B0(n42), .B1(K_r11[13]), .Y(
        K13[4]) );
  AO22X1 U1047 ( .A0(n66), .A1(K_r10[27]), .B0(K_r10[4]), .B1(n246), .Y(K12[4]) );
  AO22X1 U1048 ( .A0(n186), .A1(K_r9[47]), .B0(n112), .B1(K_r9[41]), .Y(K11[4]) );
  AO22X1 U1049 ( .A0(n172), .A1(K_r8[33]), .B0(n67), .B1(K_r8[55]), .Y(K10[4])
         );
  AO22X1 U1050 ( .A0(n77), .A1(K_r7[12]), .B0(K_r7[19]), .B1(n252), .Y(K9[4])
         );
  AO22X1 U1051 ( .A0(n196), .A1(K_r6[12]), .B0(K_r6[19]), .B1(n130), .Y(K8[4])
         );
  AO22X1 U1052 ( .A0(n148), .A1(K_r5[33]), .B0(n265), .B1(K_r5[55]), .Y(K7[4])
         );
  AO22X1 U1053 ( .A0(n38), .A1(K_r4[47]), .B0(n257), .B1(K_r4[41]), .Y(K6[4])
         );
  AO22X1 U1054 ( .A0(n159), .A1(K_r3[27]), .B0(K_r3[4]), .B1(n143), .Y(K5[4])
         );
  AO22X1 U1055 ( .A0(n68), .A1(K_r2[18]), .B0(n207), .B1(K_r2[13]), .Y(K4[4])
         );
  OAI22X1 U1056 ( .A0(n161), .A1(n400), .B0(n10), .B1(n406), .Y(K3[4]) );
  AO22X1 U1057 ( .A0(n190), .A1(K_r0[10]), .B0(n106), .B1(K_r0[46]), .Y(K2[4])
         );
  AO22X1 U1058 ( .A0(K[53]), .A1(n26), .B0(K[3]), .B1(n171), .Y(K1[4]) );
  AO22X1 U1059 ( .A0(n193), .A1(K_r14[27]), .B0(n118), .B1(K_r14[34]), .Y(
        K16[16]) );
  AO22X1 U1060 ( .A0(n263), .A1(K_r13[20]), .B0(n26), .B1(K_r13[41]), .Y(
        K15[16]) );
  AO22X1 U1061 ( .A0(n115), .A1(K_r12[55]), .B0(K_r12[6]), .B1(n178), .Y(
        K14[16]) );
  AO22X1 U1062 ( .A0(n178), .A1(K_r11[17]), .B0(n88), .B1(K_r11[12]), .Y(
        K13[16]) );
  AO22X1 U1063 ( .A0(n184), .A1(K_r10[3]), .B0(n32), .B1(K_r10[26]), .Y(
        K12[16]) );
  AO22X1 U1064 ( .A0(n87), .A1(K_r9[40]), .B0(n260), .B1(K_r9[46]), .Y(K11[16]) );
  AO22X1 U1065 ( .A0(K_r8[54]), .A1(n33), .B0(K_r8[32]), .B1(n163), .Y(K10[16]) );
  AO22X1 U1066 ( .A0(n91), .A1(K_r7[11]), .B0(n209), .B1(K_r7[18]), .Y(K9[16])
         );
  AO22X1 U1067 ( .A0(n199), .A1(K_r6[11]), .B0(n103), .B1(K_r6[18]), .Y(K8[16]) );
  AO22X1 U1068 ( .A0(n225), .A1(K_r5[54]), .B0(K_r5[32]), .B1(n150), .Y(K7[16]) );
  AO22X1 U1069 ( .A0(n195), .A1(K_r4[40]), .B0(n143), .B1(K_r4[46]), .Y(K6[16]) );
  AO22X1 U1070 ( .A0(n65), .A1(K_r3[3]), .B0(n234), .B1(K_r3[26]), .Y(K5[16])
         );
  AO22X1 U1071 ( .A0(n70), .A1(K_r2[17]), .B0(n209), .B1(K_r2[12]), .Y(K4[16])
         );
  AO22X1 U1072 ( .A0(n172), .A1(K_r1[55]), .B0(K_r1[6]), .B1(n131), .Y(K3[16])
         );
  AO22X1 U1073 ( .A0(n56), .A1(K_r0[20]), .B0(n211), .B1(K_r0[41]), .Y(K2[16])
         );
  AO22X1 U1074 ( .A0(n45), .A1(K[27]), .B0(n250), .B1(K[34]), .Y(K1[16]) );
  AO22X1 U1075 ( .A0(n195), .A1(K_r14[41]), .B0(n113), .B1(K_r14[48]), .Y(
        K16[10]) );
  AO22X1 U1076 ( .A0(n267), .A1(K_r13[34]), .B0(K_r13[55]), .B1(n148), .Y(
        K15[10]) );
  OAI22X1 U1077 ( .A0(n3), .A1(n411), .B0(n164), .B1(n419), .Y(K14[10]) );
  AO22X1 U1078 ( .A0(n122), .A1(K_r11[26]), .B0(n266), .B1(K_r11[6]), .Y(
        K13[10]) );
  AO22X1 U1079 ( .A0(n185), .A1(K_r10[17]), .B0(n116), .B1(K_r10[40]), .Y(
        K12[10]) );
  AO22X1 U1080 ( .A0(n173), .A1(K_r9[3]), .B0(K_r9[54]), .B1(n120), .Y(K11[10]) );
  AO22X1 U1081 ( .A0(n169), .A1(K_r8[46]), .B0(n98), .B1(K_r8[11]), .Y(K10[10]) );
  AO22X1 U1082 ( .A0(n93), .A1(K_r7[25]), .B0(n157), .B1(K_r7[32]), .Y(K9[10])
         );
  AO22X1 U1083 ( .A0(n200), .A1(K_r6[25]), .B0(n17), .B1(K_r6[32]), .Y(K8[10])
         );
  AO22X1 U1084 ( .A0(n36), .A1(K_r5[46]), .B0(n184), .B1(K_r5[11]), .Y(K7[10])
         );
  AO22X1 U1085 ( .A0(n50), .A1(K_r4[3]), .B0(K_r4[54]), .B1(n259), .Y(K6[10])
         );
  AO22X1 U1086 ( .A0(n67), .A1(K_r3[17]), .B0(n220), .B1(K_r3[40]), .Y(K5[10])
         );
  AO22X1 U1087 ( .A0(n170), .A1(K_r2[26]), .B0(n113), .B1(K_r2[6]), .Y(K4[10])
         );
  OAI22X1 U1088 ( .A0(n157), .A1(n410), .B0(n18), .B1(n418), .Y(K3[10]) );
  AO22X1 U1089 ( .A0(n55), .A1(K_r0[34]), .B0(K_r0[55]), .B1(n205), .Y(K2[10])
         );
  AO22X1 U1090 ( .A0(n44), .A1(K[41]), .B0(n200), .B1(K[48]), .Y(K1[10]) );
  AO22X1 U1091 ( .A0(n94), .A1(K_r14[24]), .B0(n180), .B1(K_r14[17]), .Y(
        K16[21]) );
  AO22X1 U1092 ( .A0(n74), .A1(K_r13[6]), .B0(n247), .B1(K_r13[10]), .Y(
        K15[21]) );
  OAI22X1 U1093 ( .A0(decrypt), .A1(n381), .B0(n167), .B1(n411), .Y(K14[21])
         );
  AO22X1 U1094 ( .A0(n108), .A1(K_r11[34]), .B0(n254), .B1(K_r11[39]), .Y(
        K13[21]) );
  AO22X1 U1095 ( .A0(n99), .A1(K_r10[48]), .B0(n252), .B1(K_r10[25]), .Y(
        K12[21]) );
  AO22X1 U1096 ( .A0(n190), .A1(K_r9[11]), .B0(K_r9[5]), .B1(n120), .Y(K11[21]) );
  AO22X1 U1097 ( .A0(n168), .A1(K_r8[54]), .B0(K_r8[19]), .B1(n132), .Y(
        K10[21]) );
  AO22X1 U1098 ( .A0(n194), .A1(K_r7[40]), .B0(n128), .B1(K_r7[33]), .Y(K9[21]) );
  AO22X1 U1099 ( .A0(n86), .A1(K_r6[40]), .B0(n225), .B1(K_r6[33]), .Y(K8[21])
         );
  AO22X1 U1100 ( .A0(K_r5[54]), .A1(n90), .B0(K_r5[19]), .B1(n265), .Y(K7[21])
         );
  AO22X1 U1101 ( .A0(n45), .A1(K_r4[11]), .B0(K_r4[5]), .B1(n258), .Y(K6[21])
         );
  AO22X1 U1102 ( .A0(n216), .A1(K_r3[48]), .B0(n59), .B1(K_r3[25]), .Y(K5[21])
         );
  AO22X1 U1103 ( .A0(n171), .A1(K_r2[34]), .B0(n115), .B1(K_r2[39]), .Y(K4[21]) );
  OAI22X1 U1104 ( .A0(n159), .A1(n380), .B0(n13), .B1(n410), .Y(K3[21]) );
  AO22X1 U1105 ( .A0(n182), .A1(K_r0[6]), .B0(n105), .B1(K_r0[10]), .Y(K2[21])
         );
  AO22X1 U1106 ( .A0(n173), .A1(K[24]), .B0(n115), .B1(K[17]), .Y(K1[21]) );
  AO22X1 U1107 ( .A0(n205), .A1(K_r14[47]), .B0(n116), .B1(K_r14[54]), .Y(
        K16[9]) );
  AO22X1 U1108 ( .A0(n195), .A1(K_r13[40]), .B0(K_r13[4]), .B1(n152), .Y(
        K15[9]) );
  AO22X1 U1109 ( .A0(n193), .A1(K_r12[26]), .B0(K_r12[18]), .B1(n147), .Y(
        K14[9]) );
  AO22X1 U1110 ( .A0(n183), .A1(K_r11[12]), .B0(n36), .B1(K_r11[32]), .Y(
        K13[9]) );
  AO22X1 U1111 ( .A0(n151), .A1(K_r10[46]), .B0(n270), .B1(K_r10[55]), .Y(
        K12[9]) );
  AO22X1 U1112 ( .A0(n185), .A1(K_r9[41]), .B0(n31), .B1(K_r9[3]), .Y(K11[9])
         );
  AO22X1 U1113 ( .A0(n84), .A1(K_r8[17]), .B0(n214), .B1(K_r8[27]), .Y(K10[9])
         );
  AO22X1 U1114 ( .A0(K_r7[6]), .A1(n23), .B0(n272), .B1(K_r7[13]), .Y(K9[9])
         );
  AO22X1 U1115 ( .A0(n195), .A1(K_r6[6]), .B0(n122), .B1(K_r6[13]), .Y(K8[9])
         );
  AO22X1 U1116 ( .A0(n200), .A1(K_r5[17]), .B0(n104), .B1(K_r5[27]), .Y(K7[9])
         );
  AO22X1 U1117 ( .A0(n65), .A1(K_r4[41]), .B0(n265), .B1(K_r4[3]), .Y(K6[9])
         );
  AO22X1 U1118 ( .A0(n158), .A1(K_r3[46]), .B0(n87), .B1(K_r3[55]), .Y(K5[9])
         );
  AO22X1 U1119 ( .A0(n67), .A1(K_r2[12]), .B0(n207), .B1(K_r2[32]), .Y(K4[9])
         );
  AO22X1 U1120 ( .A0(K_r1[26]), .A1(n34), .B0(K_r1[18]), .B1(n249), .Y(K3[9])
         );
  AO22X1 U1121 ( .A0(n65), .A1(K_r0[40]), .B0(K_r0[4]), .B1(n252), .Y(K2[9])
         );
  AO22X1 U1122 ( .A0(n54), .A1(K[47]), .B0(n212), .B1(K[54]), .Y(K1[9]) );
  AO22X1 U1123 ( .A0(n49), .A1(K_r14[26]), .B0(n249), .B1(K_r14[19]), .Y(
        K16[3]) );
  AO22X1 U1124 ( .A0(n38), .A1(K_r13[33]), .B0(n266), .B1(K_r13[12]), .Y(
        K15[3]) );
  AO22X1 U1125 ( .A0(n236), .A1(K_r12[55]), .B0(K_r12[47]), .B1(n146), .Y(
        K14[3]) );
  AO22X1 U1126 ( .A0(n182), .A1(K_r11[41]), .B0(K_r11[4]), .B1(n142), .Y(
        K13[3]) );
  AO22X1 U1127 ( .A0(n50), .A1(K_r10[18]), .B0(n268), .B1(K_r10[27]), .Y(
        K12[3]) );
  AO22X1 U1128 ( .A0(n187), .A1(K_r9[13]), .B0(n128), .B1(K_r9[32]), .Y(K11[3]) );
  AO22X1 U1129 ( .A0(n231), .A1(K_r8[24]), .B0(n22), .B1(K_r8[46]), .Y(K10[3])
         );
  AO22X1 U1130 ( .A0(n191), .A1(K_r7[10]), .B0(n79), .B1(K_r7[3]), .Y(K9[3])
         );
  AO22X1 U1131 ( .A0(n97), .A1(K_r6[10]), .B0(n207), .B1(K_r6[3]), .Y(K8[3])
         );
  AO22X1 U1132 ( .A0(n202), .A1(K_r5[46]), .B0(n1), .B1(K_r5[24]), .Y(K7[3])
         );
  AO22X1 U1133 ( .A0(n171), .A1(K_r4[32]), .B0(n48), .B1(K_r4[13]), .Y(K6[3])
         );
  AO22X1 U1134 ( .A0(n224), .A1(K_r3[18]), .B0(n106), .B1(K_r3[27]), .Y(K5[3])
         );
  AO22X1 U1135 ( .A0(n71), .A1(K_r2[41]), .B0(K_r2[4]), .B1(n239), .Y(K4[3])
         );
  AO22X1 U1136 ( .A0(K_r1[55]), .A1(n33), .B0(K_r1[47]), .B1(n158), .Y(K3[3])
         );
  AO22X1 U1137 ( .A0(n187), .A1(K_r0[33]), .B0(n103), .B1(K_r0[12]), .Y(K2[3])
         );
  AO22X1 U1138 ( .A0(n177), .A1(K[26]), .B0(n110), .B1(K[19]), .Y(K1[3]) );
  AO22X1 U1139 ( .A0(n200), .A1(K_r14[35]), .B0(K_r14[42]), .B1(n156), .Y(
        K16[41]) );
  AO22X1 U1140 ( .A0(n199), .A1(K_r13[28]), .B0(n115), .B1(K_r13[49]), .Y(
        K15[41]) );
  OAI22X1 U1141 ( .A0(n161), .A1(n423), .B0(n17), .B1(n415), .Y(K14[41]) );
  AO22X1 U1142 ( .A0(n111), .A1(K_r11[22]), .B0(n242), .B1(K_r11[0]), .Y(
        K13[41]) );
  AO22X1 U1143 ( .A0(n181), .A1(K_r10[45]), .B0(n61), .B1(K_r10[36]), .Y(
        K12[41]) );
  AO22X1 U1144 ( .A0(K_r9[50]), .A1(n28), .B0(K_r9[31]), .B1(n241), .Y(K11[41]) );
  AO22X1 U1145 ( .A0(n82), .A1(K_r8[9]), .B0(n214), .B1(K_r8[44]), .Y(K10[41])
         );
  AO22X1 U1146 ( .A0(n79), .A1(K_r7[23]), .B0(K_r7[30]), .B1(n179), .Y(K9[41])
         );
  AO22X1 U1147 ( .A0(n196), .A1(K_r6[23]), .B0(K_r6[30]), .B1(n131), .Y(K8[41]) );
  AO22X1 U1148 ( .A0(n202), .A1(K_r5[9]), .B0(n156), .B1(K_r5[44]), .Y(K7[41])
         );
  AO22X1 U1149 ( .A0(n228), .A1(K_r4[50]), .B0(K_r4[31]), .B1(n155), .Y(K6[41]) );
  AO22X1 U1150 ( .A0(n54), .A1(K_r3[45]), .B0(n206), .B1(K_r3[36]), .Y(K5[41])
         );
  AO22X1 U1151 ( .A0(n167), .A1(K_r2[22]), .B0(n20), .B1(K_r2[0]), .Y(K4[41])
         );
  OAI22X1 U1152 ( .A0(n5), .A1(n422), .B0(n165), .B1(n414), .Y(K3[41]) );
  AO22X1 U1153 ( .A0(n62), .A1(K_r0[28]), .B0(n210), .B1(K_r0[49]), .Y(K2[41])
         );
  AO22X1 U1154 ( .A0(n51), .A1(K[35]), .B0(K[42]), .B1(n185), .Y(K1[41]) );
  AO22X1 U1155 ( .A0(n193), .A1(K_r14[51]), .B0(n112), .B1(K_r14[31]), .Y(
        K16[26]) );
  AO22X1 U1156 ( .A0(n41), .A1(K_r13[38]), .B0(n246), .B1(K_r13[44]), .Y(
        K15[26]) );
  AO22X1 U1157 ( .A0(n136), .A1(K_r12[52]), .B0(n264), .B1(K_r12[30]), .Y(
        K14[26]) );
  AO22X1 U1158 ( .A0(n177), .A1(K_r11[16]), .B0(K_r11[7]), .B1(n140), .Y(
        K13[26]) );
  AO22X1 U1159 ( .A0(n183), .A1(K_r10[2]), .B0(n54), .B1(K_r10[21]), .Y(
        K12[26]) );
  AO22X1 U1160 ( .A0(n189), .A1(K_r9[43]), .B0(K_r9[35]), .B1(n123), .Y(
        K11[26]) );
  AO22X1 U1161 ( .A0(n78), .A1(K_r8[49]), .B0(n213), .B1(K_r8[29]), .Y(K10[26]) );
  AO22X1 U1162 ( .A0(n86), .A1(K_r7[8]), .B0(n256), .B1(K_r7[15]), .Y(K9[26])
         );
  AO22X1 U1163 ( .A0(n198), .A1(K_r6[8]), .B0(n13), .B1(K_r6[15]), .Y(K8[26])
         );
  AO22X1 U1164 ( .A0(n203), .A1(K_r5[49]), .B0(n88), .B1(K_r5[29]), .Y(K7[26])
         );
  AO22X1 U1165 ( .A0(K_r4[43]), .A1(n22), .B0(K_r4[35]), .B1(n159), .Y(K6[26])
         );
  AO22X1 U1166 ( .A0(n61), .A1(K_r3[2]), .B0(n206), .B1(K_r3[21]), .Y(K5[26])
         );
  AO22X1 U1167 ( .A0(n73), .A1(K_r2[16]), .B0(K_r2[7]), .B1(n167), .Y(K4[26])
         );
  AO22X1 U1168 ( .A0(n171), .A1(K_r1[52]), .B0(n110), .B1(K_r1[30]), .Y(K3[26]) );
  AO22X1 U1169 ( .A0(n183), .A1(K_r0[38]), .B0(n104), .B1(K_r0[44]), .Y(K2[26]) );
  AO22X1 U1170 ( .A0(n48), .A1(K[51]), .B0(n268), .B1(K[31]), .Y(K1[26]) );
  AO22X1 U1171 ( .A0(n42), .A1(K_r14[7]), .B0(n259), .B1(K_r14[0]), .Y(K16[47]) );
  AO22X1 U1172 ( .A0(n36), .A1(K_r13[14]), .B0(K_r13[52]), .B1(n200), .Y(
        K15[47]) );
  AO22X1 U1173 ( .A0(n141), .A1(K_r12[28]), .B0(n268), .B1(K_r12[38]), .Y(
        K14[47]) );
  AO22X1 U1174 ( .A0(n140), .A1(K_r11[42]), .B0(n255), .B1(K_r11[51]), .Y(
        K13[47]) );
  AO22X1 U1175 ( .A0(n89), .A1(K_r10[1]), .B0(n260), .B1(K_r10[37]), .Y(
        K12[47]) );
  AO22X1 U1176 ( .A0(n95), .A1(K_r9[15]), .B0(K_r9[23]), .B1(n262), .Y(K11[47]) );
  AO22X1 U1177 ( .A0(n83), .A1(K_r8[29]), .B0(n214), .B1(K_r8[9]), .Y(K10[47])
         );
  AO22X1 U1178 ( .A0(n190), .A1(K_r7[50]), .B0(n146), .B1(K_r7[43]), .Y(K9[47]) );
  AO22X1 U1179 ( .A0(n96), .A1(K_r6[50]), .B0(n258), .B1(K_r6[43]), .Y(K8[47])
         );
  AO22X1 U1180 ( .A0(n201), .A1(K_r5[29]), .B0(n150), .B1(K_r5[9]), .Y(K7[47])
         );
  AO22X1 U1181 ( .A0(n204), .A1(K_r4[15]), .B0(K_r4[23]), .B1(n153), .Y(K6[47]) );
  AO22X1 U1182 ( .A0(n223), .A1(K_r3[1]), .B0(n55), .B1(K_r3[37]), .Y(K5[47])
         );
  AO22X1 U1183 ( .A0(n165), .A1(K_r2[42]), .B0(n8), .B1(K_r2[51]), .Y(K4[47])
         );
  AO22X1 U1184 ( .A0(n69), .A1(K_r1[38]), .B0(n209), .B1(K_r1[28]), .Y(K3[47])
         );
  AO22X1 U1185 ( .A0(n189), .A1(K_r0[14]), .B0(K_r0[52]), .B1(n128), .Y(K2[47]) );
  AO22X1 U1186 ( .A0(n178), .A1(K[7]), .B0(n108), .B1(K[0]), .Y(K1[47]) );
  AO22X1 U1187 ( .A0(n194), .A1(K_r14[1]), .B0(K_r14[8]), .B1(n155), .Y(
        K16[28]) );
  AO22X1 U1188 ( .A0(n203), .A1(K_r13[49]), .B0(n70), .B1(K_r13[15]), .Y(
        K15[28]) );
  OAI22X1 U1189 ( .A0(n1), .A1(n399), .B0(n167), .B1(n403), .Y(K14[28]) );
  AO22X1 U1190 ( .A0(K_r11[43]), .A1(n19), .B0(K_r11[21]), .B1(n193), .Y(
        K13[28]) );
  AO22X1 U1191 ( .A0(n38), .A1(K_r10[2]), .B0(n263), .B1(K_r10[7]), .Y(K12[28]) );
  AO22X1 U1192 ( .A0(n189), .A1(K_r9[52]), .B0(n63), .B1(K_r9[16]), .Y(K11[28]) );
  AO22X1 U1193 ( .A0(n170), .A1(K_r8[38]), .B0(n84), .B1(K_r8[30]), .Y(K10[28]) );
  AO22X1 U1194 ( .A0(n85), .A1(K_r7[44]), .B0(K_r7[51]), .B1(n241), .Y(K9[28])
         );
  AO22X1 U1195 ( .A0(n198), .A1(K_r6[44]), .B0(K_r6[51]), .B1(n137), .Y(K8[28]) );
  AO22X1 U1196 ( .A0(n34), .A1(K_r5[38]), .B0(n270), .B1(K_r5[30]), .Y(K7[28])
         );
  AO22X1 U1197 ( .A0(n42), .A1(K_r4[52]), .B0(n204), .B1(K_r4[16]), .Y(K6[28])
         );
  AO22X1 U1198 ( .A0(n224), .A1(K_r3[2]), .B0(n154), .B1(K_r3[7]), .Y(K5[28])
         );
  AO22X1 U1199 ( .A0(n173), .A1(K_r2[43]), .B0(K_r2[21]), .B1(n134), .Y(K4[28]) );
  OAI22X1 U1200 ( .A0(n160), .A1(n398), .B0(n16), .B1(n402), .Y(K3[28]) );
  AO22X1 U1201 ( .A0(n59), .A1(K_r0[49]), .B0(n210), .B1(K_r0[15]), .Y(K2[28])
         );
  AO22X1 U1202 ( .A0(n49), .A1(K[1]), .B0(K[8]), .B1(n179), .Y(K1[28]) );
  CLKINVX1 U1203 ( .A(decrypt), .Y(n272) );
endmodule


module sbox1_0 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n69, n70, n71,
         n72;

  OAI222X4 U13 ( .A0(addr[5]), .A1(n40), .B0(n1), .B1(n41), .C0(n42), .C1(n72), 
        .Y(dout[3]) );
  OAI21X2 U42 ( .A0(n4), .A1(n29), .B0(n35), .Y(n18) );
  NAND2X2 U44 ( .A(addr[6]), .B(n9), .Y(n26) );
  NAND2X2 U48 ( .A(addr[1]), .B(n12), .Y(n27) );
  OAI22X2 U49 ( .A0(n6), .A1(n71), .B0(addr[5]), .B1(n21), .Y(n56) );
  NAND2X2 U50 ( .A(n3), .B(n6), .Y(n21) );
  NOR2X2 U51 ( .A(n6), .B(n3), .Y(n17) );
  NOR3X2 U55 ( .A(n2), .B(addr[6]), .C(n72), .Y(n39) );
  NOR2X2 U56 ( .A(n32), .B(n3), .Y(n48) );
  NAND2X2 U57 ( .A(addr[1]), .B(addr[6]), .Y(n32) );
  NAND2X2 U59 ( .A(n9), .B(n12), .Y(n29) );
  NOR2X1 U1 ( .A(n27), .B(n21), .Y(n37) );
  BUFX4 U2 ( .A(addr[4]), .Y(n2) );
  CLKBUFX3 U3 ( .A(addr[2]), .Y(n1) );
  OAI32X1 U4 ( .A0(n29), .A1(n2), .A2(n4), .B0(n26), .B1(n28), .Y(n61) );
  NOR2BXL U5 ( .AN(n23), .B(n1), .Y(n19) );
  CLKBUFX3 U6 ( .A(addr[2]), .Y(n4) );
  INVX3 U7 ( .A(addr[6]), .Y(n12) );
  OAI221X4 U8 ( .A0(n53), .A1(n71), .B0(addr[5]), .B1(n54), .C0(n55), .Y(
        dout[2]) );
  OAI221X4 U9 ( .A0(addr[5]), .A1(n14), .B0(n15), .B1(n71), .C0(n16), .Y(
        dout[4]) );
  OA21XL U10 ( .A0(n46), .A1(n26), .B0(n34), .Y(n22) );
  AOI222XL U11 ( .A0(n8), .A1(n1), .B0(n2), .B1(n31), .C0(n10), .C1(n72), .Y(
        n30) );
  AOI2BB2X1 U12 ( .B0(n2), .B1(n10), .A0N(addr[4]), .A1N(n26), .Y(n50) );
  BUFX4 U14 ( .A(addr[3]), .Y(n3) );
  CLKINVX1 U15 ( .A(n29), .Y(n8) );
  CLKINVX1 U16 ( .A(n28), .Y(n13) );
  NAND2BX1 U17 ( .AN(n37), .B(n22), .Y(n57) );
  CLKXOR2X2 U18 ( .A(n69), .B(n72), .Y(n51) );
  NOR2X1 U19 ( .A(n6), .B(n69), .Y(n23) );
  OAI21XL U20 ( .A0(n69), .A1(n27), .B0(n50), .Y(n49) );
  NAND2X1 U21 ( .A(n48), .B(n6), .Y(n34) );
  NAND2X1 U22 ( .A(n72), .B(n69), .Y(n28) );
  OAI211X1 U23 ( .A0(n6), .A1(n27), .B0(n33), .C0(n34), .Y(n52) );
  CLKINVX1 U24 ( .A(n32), .Y(n10) );
  NAND2X1 U25 ( .A(n17), .B(n7), .Y(n33) );
  CLKINVX1 U26 ( .A(n27), .Y(n11) );
  CLKINVX1 U27 ( .A(n26), .Y(n7) );
  CLKINVX1 U28 ( .A(n46), .Y(n70) );
  AO22X1 U29 ( .A0(n51), .A1(n7), .B0(n69), .B1(n18), .Y(n65) );
  OAI31X1 U30 ( .A0(n72), .A1(n3), .A2(n9), .B0(n38), .Y(n36) );
  AOI31XL U31 ( .A0(n9), .A1(n72), .A2(n2), .B0(n39), .Y(n38) );
  AOI211X1 U32 ( .A0(n5), .A1(n4), .B0(n24), .C0(n25), .Y(n15) );
  CLKINVX1 U33 ( .A(n33), .Y(n5) );
  AOI211X1 U34 ( .A0(n26), .A1(n27), .B0(n28), .C0(n2), .Y(n25) );
  OAI22X1 U35 ( .A0(n21), .A1(n29), .B0(n30), .B1(n69), .Y(n24) );
  AOI211X1 U36 ( .A0(n10), .A1(n23), .B0(n60), .C0(n61), .Y(n53) );
  OAI22X1 U37 ( .A0(n50), .A1(n72), .B0(n3), .B1(n35), .Y(n60) );
  CLKINVX3 U38 ( .A(addr[5]), .Y(n71) );
  NAND2X1 U39 ( .A(n3), .B(n71), .Y(n46) );
  NAND2X1 U40 ( .A(n11), .B(n1), .Y(n35) );
  XOR2X1 U41 ( .A(n59), .B(n2), .Y(n58) );
  NAND2X1 U43 ( .A(n1), .B(n3), .Y(n59) );
  OAI22XL U45 ( .A0(n3), .A1(n9), .B0(n69), .B1(n29), .Y(n47) );
  AOI211XL U46 ( .A0(n43), .A1(n69), .B0(n44), .C0(n37), .Y(n42) );
  OAI22XL U47 ( .A0(n45), .A1(n6), .B0(n46), .B1(n32), .Y(n44) );
  OAI22XL U52 ( .A0(n12), .A1(n71), .B0(n2), .B1(addr[1]), .Y(n43) );
  AOI221XL U53 ( .A0(n70), .A1(addr[6]), .B0(addr[5]), .B1(n47), .C0(n48), .Y(
        n45) );
  OAI21XL U54 ( .A0(addr[1]), .A1(n21), .B0(n22), .Y(n20) );
  AOI221XL U58 ( .A0(n8), .A1(n23), .B0(n48), .B1(n71), .C0(n66), .Y(n63) );
  OAI31X1 U60 ( .A0(n71), .A1(n2), .A2(n67), .B0(n68), .Y(n66) );
  OA21XL U61 ( .A0(n3), .A1(n12), .B0(n32), .Y(n67) );
  OAI21XL U62 ( .A0(n17), .A1(n56), .B0(n11), .Y(n68) );
  OAI21XL U63 ( .A0(n1), .A1(n9), .B0(n32), .Y(n31) );
  INVX4 U64 ( .A(n4), .Y(n72) );
  AOI222XL U65 ( .A0(n17), .A1(n18), .B0(n19), .B1(addr[6]), .C0(n1), .C1(n20), 
        .Y(n16) );
  NOR4BBX1 U66 ( .AN(n34), .BN(n35), .C(n36), .D(n37), .Y(n14) );
  AOI222XL U67 ( .A0(n8), .A1(n51), .B0(n52), .B1(n72), .C0(n18), .C1(n6), .Y(
        n40) );
  AOI2BB2XL U68 ( .B0(addr[5]), .B1(n49), .A0N(n21), .A1N(addr[1]), .Y(n41) );
  AOI32X1 U69 ( .A0(n4), .A1(n56), .A2(n8), .B0(n57), .B1(n72), .Y(n55) );
  AOI222XL U70 ( .A0(n17), .A1(n9), .B0(n58), .B1(addr[1]), .C0(n13), .C1(n12), 
        .Y(n54) );
  OAI221X1 U71 ( .A0(n62), .A1(n71), .B0(n4), .B1(n63), .C0(n64), .Y(dout[1])
         );
  AOI32XL U72 ( .A0(addr[6]), .A1(n56), .A2(n1), .B0(n65), .B1(n71), .Y(n64)
         );
  AOI221X1 U73 ( .A0(n8), .A1(n51), .B0(n4), .B1(n48), .C0(n39), .Y(n62) );
  CLKINVX3 U74 ( .A(n2), .Y(n6) );
  CLKINVX3 U75 ( .A(addr[1]), .Y(n9) );
  CLKINVX3 U76 ( .A(n3), .Y(n69) );
endmodule


module sbox2_0 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n81, n82, n83;

  NAND2X2 U55 ( .A(n2), .B(n6), .Y(n28) );
  NAND2X2 U57 ( .A(addr[2]), .B(n11), .Y(n60) );
  NAND2X2 U60 ( .A(addr[5]), .B(addr[2]), .Y(n32) );
  NOR2X2 U61 ( .A(n16), .B(n13), .Y(n63) );
  NAND2X2 U62 ( .A(n15), .B(n83), .Y(n18) );
  NAND2X2 U63 ( .A(n3), .B(n82), .Y(n40) );
  NAND2X2 U64 ( .A(addr[6]), .B(n15), .Y(n42) );
  NAND2X2 U67 ( .A(n3), .B(n2), .Y(n31) );
  AOI222XL U1 ( .A0(n5), .A1(n81), .B0(n76), .B1(n82), .C0(n24), .C1(n13), .Y(
        n75) );
  CLKINVX1 U2 ( .A(n43), .Y(n16) );
  AOI211X1 U3 ( .A0(n12), .A1(n69), .B0(n70), .C0(n71), .Y(n68) );
  NOR2X1 U4 ( .A(n60), .B(n2), .Y(n23) );
  NOR2X1 U5 ( .A(n40), .B(n2), .Y(n24) );
  CLKBUFX4 U6 ( .A(addr[4]), .Y(n2) );
  CLKINVX1 U7 ( .A(addr[5]), .Y(n1) );
  OAI22X1 U8 ( .A0(n47), .A1(n50), .B0(n75), .B1(n11), .Y(n70) );
  INVX3 U9 ( .A(addr[5]), .Y(n11) );
  OAI211X4 U10 ( .A0(n17), .A1(n18), .B0(n19), .C0(n20), .Y(dout[4]) );
  NAND2X1 U11 ( .A(addr[1]), .B(addr[6]), .Y(n43) );
  CLKINVX2 U12 ( .A(addr[1]), .Y(n15) );
  OAI221X1 U13 ( .A0(addr[1]), .A1(n28), .B0(n31), .B1(n15), .C0(n77), .Y(n69)
         );
  NAND2X4 U14 ( .A(addr[1]), .B(n83), .Y(n50) );
  INVX3 U15 ( .A(addr[6]), .Y(n83) );
  NAND2XL U16 ( .A(n62), .B(n6), .Y(n55) );
  AOI2BB2X1 U17 ( .B0(n11), .B1(n8), .A0N(n60), .A1N(n28), .Y(n47) );
  NOR3BXL U18 ( .AN(n29), .B(n30), .C(n5), .Y(n17) );
  BUFX4 U19 ( .A(addr[3]), .Y(n3) );
  NAND2X1 U20 ( .A(n5), .B(n16), .Y(n51) );
  CLKINVX1 U21 ( .A(n18), .Y(n13) );
  CLKINVX1 U22 ( .A(n49), .Y(n5) );
  CLKINVX1 U23 ( .A(n42), .Y(n14) );
  OAI31X1 U24 ( .A0(n40), .A1(n83), .A2(n11), .B0(n41), .Y(n36) );
  OAI21XL U25 ( .A0(n1), .A1(n15), .B0(n24), .Y(n41) );
  OAI22X1 U26 ( .A0(n42), .A1(n40), .B0(n63), .B1(n32), .Y(n80) );
  INVX1 U27 ( .A(n50), .Y(n81) );
  OAI22X1 U28 ( .A0(n42), .A1(n6), .B0(n9), .B1(n43), .Y(n35) );
  NAND3X1 U29 ( .A(n9), .B(n11), .C(n15), .Y(n53) );
  NAND2X1 U30 ( .A(n6), .B(n9), .Y(n49) );
  OAI21XL U31 ( .A0(n82), .A1(n31), .B0(n29), .Y(n79) );
  OAI22XL U32 ( .A0(n47), .A1(n18), .B0(n48), .B1(n32), .Y(n46) );
  AOI222XL U33 ( .A0(n81), .A1(n49), .B0(n7), .B1(n83), .C0(n5), .C1(n13), .Y(
        n48) );
  CLKINVX1 U34 ( .A(n60), .Y(n10) );
  OAI2BB2XL U35 ( .B0(n50), .B1(n29), .A0N(n38), .A1N(n7), .Y(n58) );
  OAI21XL U36 ( .A0(n52), .A1(n50), .B0(n53), .Y(n44) );
  OAI21XL U37 ( .A0(n31), .A1(n50), .B0(n51), .Y(n45) );
  CLKINVX1 U38 ( .A(n40), .Y(n8) );
  CLKINVX1 U39 ( .A(n28), .Y(n4) );
  CLKINVX1 U40 ( .A(n31), .Y(n7) );
  CLKINVX1 U41 ( .A(n32), .Y(n12) );
  AOI2BB1X1 U42 ( .A0N(n38), .A1N(n39), .B0(n28), .Y(n37) );
  OAI22XL U43 ( .A0(n60), .A1(n50), .B0(n63), .B1(n32), .Y(n62) );
  AO21XL U44 ( .A0(n82), .A1(n4), .B0(n23), .Y(n78) );
  AO21X1 U45 ( .A0(n6), .A1(n10), .B0(n24), .Y(n22) );
  NAND3X1 U46 ( .A(n82), .B(n9), .C(addr[5]), .Y(n29) );
  OAI22X1 U47 ( .A0(addr[5]), .A1(n43), .B0(n42), .B1(n11), .Y(n38) );
  AOI2BB1X1 U48 ( .A0N(n3), .A1N(n1), .B0(n4), .Y(n52) );
  NOR3X1 U49 ( .A(addr[1]), .B(addr[2]), .C(n11), .Y(n39) );
  AOI2BB1XL U50 ( .A0N(n72), .A1N(n73), .B0(addr[5]), .Y(n71) );
  OAI31XL U51 ( .A0(n50), .A1(n2), .A2(n6), .B0(n74), .Y(n73) );
  OAI21XL U52 ( .A0(n7), .A1(n8), .B0(n14), .Y(n74) );
  NAND2X1 U53 ( .A(n81), .B(n2), .Y(n27) );
  OAI31XL U54 ( .A0(n63), .A1(n3), .A2(addr[2]), .B0(n51), .Y(n72) );
  OAI211X1 U56 ( .A0(n25), .A1(n11), .B0(n26), .C0(n27), .Y(n21) );
  NAND3X1 U58 ( .A(n9), .B(n11), .C(addr[6]), .Y(n26) );
  AOI2BB2X1 U59 ( .B0(n14), .B1(n6), .A0N(n15), .A1N(n28), .Y(n25) );
  OAI22XL U65 ( .A0(addr[5]), .A1(n31), .B0(n3), .B1(n32), .Y(n30) );
  OAI2BB2XL U66 ( .B0(n52), .B1(n42), .A0N(n1), .A1N(n65), .Y(n64) );
  OAI211X1 U68 ( .A0(n18), .A1(n2), .B0(n27), .C0(n51), .Y(n65) );
  NAND3X1 U69 ( .A(n14), .B(n9), .C(n3), .Y(n77) );
  AOI2BB2XL U70 ( .B0(n3), .B1(n59), .A0N(n27), .A1N(n32), .Y(n56) );
  OAI211XL U71 ( .A0(n60), .A1(n18), .B0(n61), .C0(n53), .Y(n59) );
  NAND3XL U72 ( .A(addr[5]), .B(n9), .C(n16), .Y(n61) );
  OAI22XL U73 ( .A0(n3), .A1(n50), .B0(n83), .B1(n49), .Y(n76) );
  NAND4X1 U74 ( .A(n54), .B(n55), .C(n56), .D(n57), .Y(dout[2]) );
  AOI32XL U75 ( .A0(addr[1]), .A1(addr[2]), .A2(n4), .B0(n64), .B1(n82), .Y(
        n54) );
  AOI221XL U76 ( .A0(n39), .A1(addr[4]), .B0(n23), .B1(n14), .C0(n58), .Y(n57)
         );
  AOI33XL U77 ( .A0(n14), .A1(n10), .A2(n2), .B0(n12), .B1(n18), .B2(n3), .Y(
        n19) );
  AOI222XL U78 ( .A0(n21), .A1(n82), .B0(n16), .B1(n22), .C0(n81), .C1(n23), 
        .Y(n20) );
  NAND3X1 U79 ( .A(n66), .B(n67), .C(n68), .Y(dout[1]) );
  AOI32XL U80 ( .A0(n10), .A1(n15), .A2(n5), .B0(n13), .B1(n78), .Y(n67) );
  AOI22X1 U81 ( .A0(n16), .A1(n79), .B0(n2), .B1(n80), .Y(n66) );
  NAND2X1 U82 ( .A(n33), .B(n34), .Y(dout[3]) );
  AOI221XL U83 ( .A0(n44), .A1(n82), .B0(addr[2]), .B1(n45), .C0(n46), .Y(n33)
         );
  AOI211X1 U84 ( .A0(n10), .A1(n35), .B0(n36), .C0(n37), .Y(n34) );
  CLKINVX3 U85 ( .A(n3), .Y(n6) );
  CLKINVX3 U86 ( .A(n2), .Y(n9) );
  CLKINVX3 U87 ( .A(addr[2]), .Y(n82) );
endmodule


module sbox3_0 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n76, n77, n78;

  NOR2X2 U35 ( .A(n16), .B(addr[3]), .Y(n46) );
  NOR2X2 U50 ( .A(addr[1]), .B(addr[6]), .Y(n47) );
  NOR2X2 U52 ( .A(n76), .B(n2), .Y(n67) );
  NOR2X2 U56 ( .A(n76), .B(n77), .Y(n60) );
  NOR2X1 U1 ( .A(n16), .B(n76), .Y(n48) );
  OAI221X1 U2 ( .A0(n30), .A1(n16), .B0(n3), .B1(addr[1]), .C0(n13), .Y(n50)
         );
  OAI22XL U3 ( .A0(n2), .A1(n77), .B0(n3), .B1(n15), .Y(n31) );
  BUFX4 U4 ( .A(addr[4]), .Y(n2) );
  CLKBUFX3 U5 ( .A(n77), .Y(n1) );
  OAI33X1 U6 ( .A0(n18), .A1(n29), .A2(n77), .B0(n16), .B1(n60), .B2(n35), .Y(
        n75) );
  INVX3 U7 ( .A(n3), .Y(n77) );
  NOR2X1 U8 ( .A(n9), .B(n3), .Y(n63) );
  NOR2X1 U9 ( .A(n18), .B(n3), .Y(n33) );
  NOR2X1 U10 ( .A(n13), .B(n3), .Y(n59) );
  NOR2X1 U11 ( .A(n3), .B(n2), .Y(n44) );
  CLKBUFX4 U12 ( .A(addr[2]), .Y(n3) );
  OAI221X1 U13 ( .A0(addr[5]), .A1(n64), .B0(n65), .B1(n78), .C0(n66), .Y(
        dout[1]) );
  NOR2X4 U14 ( .A(n10), .B(n14), .Y(n30) );
  NOR2X4 U15 ( .A(addr[3]), .B(n2), .Y(n24) );
  NOR2X4 U16 ( .A(n14), .B(addr[6]), .Y(n29) );
  INVX3 U17 ( .A(addr[1]), .Y(n14) );
  NAND2XL U18 ( .A(n60), .B(n30), .Y(n22) );
  OAI211XL U19 ( .A0(n2), .A1(n8), .B0(n26), .C0(n27), .Y(n25) );
  NAND4XL U20 ( .A(n40), .B(n41), .C(n42), .D(n43), .Y(n39) );
  CLKINVX1 U21 ( .A(n22), .Y(n6) );
  INVX1 U22 ( .A(n30), .Y(n4) );
  CLKINVX1 U23 ( .A(n48), .Y(n15) );
  NAND2X1 U24 ( .A(n9), .B(n11), .Y(n32) );
  CLKINVX1 U25 ( .A(n68), .Y(n11) );
  CLKINVX1 U26 ( .A(n34), .Y(n20) );
  CLKINVX1 U27 ( .A(n35), .Y(n5) );
  CLKINVX1 U28 ( .A(n40), .Y(n7) );
  CLKINVX1 U29 ( .A(n47), .Y(n13) );
  NOR2X1 U30 ( .A(n9), .B(n77), .Y(n51) );
  NOR2X1 U31 ( .A(n4), .B(n77), .Y(n45) );
  INVX1 U32 ( .A(n29), .Y(n12) );
  AOI21X1 U33 ( .A0(n76), .A1(n77), .B0(n60), .Y(n34) );
  OAI21XL U34 ( .A0(n44), .A1(n24), .B0(n30), .Y(n72) );
  CLKINVX1 U36 ( .A(n73), .Y(n9) );
  NOR2X1 U37 ( .A(n12), .B(n16), .Y(n68) );
  NOR2X1 U38 ( .A(n30), .B(n47), .Y(n35) );
  OAI21XL U39 ( .A0(n45), .A1(n63), .B0(n24), .Y(n54) );
  NAND2X1 U40 ( .A(n51), .B(n67), .Y(n40) );
  CLKINVX1 U41 ( .A(n67), .Y(n18) );
  CLKINVX1 U42 ( .A(n63), .Y(n8) );
  CLKINVX1 U43 ( .A(n44), .Y(n19) );
  CLKINVX1 U44 ( .A(n33), .Y(n17) );
  OR2X1 U45 ( .A(n51), .B(n59), .Y(n28) );
  OAI221X1 U46 ( .A0(n12), .A1(n19), .B0(n77), .B1(n11), .C0(n61), .Y(n56) );
  AOI221XL U47 ( .A0(n59), .A1(n2), .B0(n62), .B1(n16), .C0(n6), .Y(n61) );
  OAI21XL U48 ( .A0(n1), .A1(n13), .B0(n8), .Y(n62) );
  XNOR2X1 U49 ( .A(addr[5]), .B(addr[3]), .Y(n52) );
  CLKINVX1 U51 ( .A(addr[5]), .Y(n78) );
  OAI221X1 U53 ( .A0(n13), .A1(n19), .B0(n4), .B1(n18), .C0(n49), .Y(n38) );
  AOI221XL U54 ( .A0(addr[3]), .A1(n50), .B0(n51), .B1(n24), .C0(n6), .Y(n49)
         );
  CLKINVX1 U55 ( .A(addr[6]), .Y(n10) );
  NAND3X1 U57 ( .A(n3), .B(n14), .C(n46), .Y(n41) );
  NOR2X1 U58 ( .A(n10), .B(addr[1]), .Y(n73) );
  AOI32XL U59 ( .A0(n1), .A1(n76), .A2(n30), .B0(n31), .B1(n10), .Y(n26) );
  AOI22XL U60 ( .A0(n2), .A1(n28), .B0(n29), .B1(n24), .Y(n27) );
  AOI222XL U61 ( .A0(n44), .A1(n29), .B0(n45), .B1(n76), .C0(n46), .C1(n47), 
        .Y(n43) );
  OAI211XL U62 ( .A0(n48), .A1(n24), .B0(n1), .C0(addr[6]), .Y(n42) );
  OAI21XL U63 ( .A0(n3), .A1(addr[1]), .B0(n12), .Y(n74) );
  AOI221XL U64 ( .A0(n68), .A1(n76), .B0(n67), .B1(n29), .C0(n69), .Y(n65) );
  OAI211X1 U65 ( .A0(n70), .A1(n77), .B0(n71), .C0(n72), .Y(n69) );
  AOI222XL U66 ( .A0(n73), .A1(n76), .B0(n47), .B1(n48), .C0(n24), .C1(n14), 
        .Y(n70) );
  OAI21XL U67 ( .A0(n63), .A1(n6), .B0(addr[4]), .Y(n71) );
  AOI221XL U68 ( .A0(n29), .A1(n20), .B0(addr[3]), .B1(n28), .C0(n58), .Y(n57)
         );
  OAI22X1 U69 ( .A0(n4), .A1(n17), .B0(n15), .B1(n9), .Y(n58) );
  OAI211X1 U70 ( .A0(n13), .A1(n17), .B0(n36), .C0(n37), .Y(dout[3]) );
  AOI32XL U71 ( .A0(n29), .A1(n3), .A2(n52), .B0(n46), .B1(n45), .Y(n36) );
  AOI22XL U72 ( .A0(n38), .A1(n78), .B0(addr[5]), .B1(n39), .Y(n37) );
  AOI221XL U73 ( .A0(n33), .A1(n29), .B0(n59), .B1(n46), .C0(n7), .Y(n66) );
  AOI221XL U74 ( .A0(n24), .A1(n74), .B0(n60), .B1(n32), .C0(n75), .Y(n64) );
  NAND4X1 U75 ( .A(n53), .B(n41), .C(n54), .D(n55), .Y(dout[2]) );
  NAND3XL U76 ( .A(n2), .B(n30), .C(n52), .Y(n53) );
  AOI2BB2XL U77 ( .B0(addr[5]), .B1(n56), .A0N(addr[5]), .A1N(n57), .Y(n55) );
  OAI221X1 U78 ( .A0(n21), .A1(n78), .B0(n2), .B1(n22), .C0(n23), .Y(dout[4])
         );
  AOI32XL U79 ( .A0(n24), .A1(n10), .A2(addr[2]), .B0(n25), .B1(n78), .Y(n23)
         );
  AOI222XL U80 ( .A0(n20), .A1(n32), .B0(n33), .B1(addr[1]), .C0(n34), .C1(n5), 
        .Y(n21) );
  CLKINVX3 U81 ( .A(n2), .Y(n16) );
  CLKINVX3 U82 ( .A(addr[3]), .Y(n76) );
endmodule


module sbox4_0 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n71,
         n72;

  OAI32X4 U12 ( .A0(n13), .A1(n2), .A2(addr[2]), .B0(n12), .B1(n35), .Y(n20)
         );
  OAI222X4 U20 ( .A0(addr[2]), .A1(n51), .B0(n37), .B1(n52), .C0(n53), .C1(n4), 
        .Y(dout[2]) );
  OAI222X4 U33 ( .A0(addr[4]), .A1(n37), .B0(n7), .B1(n35), .C0(n2), .C1(n25), 
        .Y(n60) );
  NAND2X2 U34 ( .A(addr[4]), .B(n2), .Y(n35) );
  NOR2X2 U43 ( .A(n71), .B(addr[4]), .Y(n30) );
  NOR2X2 U45 ( .A(n12), .B(n2), .Y(n32) );
  NAND2X2 U51 ( .A(n7), .B(n72), .Y(n25) );
  NOR2X2 U52 ( .A(n16), .B(addr[5]), .Y(n46) );
  NAND2X2 U53 ( .A(addr[6]), .B(addr[1]), .Y(n58) );
  NAND2X2 U54 ( .A(addr[1]), .B(n72), .Y(n27) );
  NOR2X2 U55 ( .A(n28), .B(n12), .Y(n22) );
  NAND2X2 U56 ( .A(n71), .B(n16), .Y(n28) );
  NAND2X2 U57 ( .A(addr[5]), .B(n16), .Y(n47) );
  NAND2X2 U58 ( .A(addr[6]), .B(n7), .Y(n37) );
  OAI222X1 U1 ( .A0(n13), .A1(n58), .B0(n46), .B1(n27), .C0(n16), .C1(n25), 
        .Y(n70) );
  CLKINVX1 U2 ( .A(n27), .Y(n10) );
  CLKINVX1 U3 ( .A(n71), .Y(n1) );
  CLKBUFX3 U4 ( .A(addr[3]), .Y(n2) );
  OAI31X4 U5 ( .A0(n25), .A1(n12), .A2(n16), .B0(n26), .Y(n24) );
  OAI221X1 U6 ( .A0(addr[2]), .A1(n63), .B0(n25), .B1(n38), .C0(n64), .Y(
        dout[1]) );
  INVX4 U7 ( .A(addr[5]), .Y(n12) );
  OAI31X1 U8 ( .A0(n35), .A1(addr[5]), .A2(n6), .B0(n36), .Y(n34) );
  AOI222XL U9 ( .A0(n16), .A1(n72), .B0(n30), .B1(n7), .C0(addr[1]), .C1(n71), 
        .Y(n29) );
  OAI222X1 U10 ( .A0(addr[1]), .A1(n59), .B0(n58), .B1(n69), .C0(n71), .C1(n36), .Y(n68) );
  NAND2XL U11 ( .A(n1), .B(addr[5]), .Y(n59) );
  AOI211XL U13 ( .A0(n60), .A1(n12), .B0(n61), .C0(n8), .Y(n51) );
  NAND2XL U14 ( .A(n16), .B(n12), .Y(n69) );
  CLKINVX1 U15 ( .A(n25), .Y(n5) );
  CLKINVX1 U16 ( .A(n28), .Y(n15) );
  CLKINVX1 U17 ( .A(n31), .Y(n3) );
  OAI21X1 U18 ( .A0(n10), .A1(n6), .B0(n4), .Y(n31) );
  AOI22X1 U19 ( .A0(n11), .A1(n32), .B0(n6), .B1(n30), .Y(n50) );
  OAI211X1 U21 ( .A0(n7), .A1(n28), .B0(n50), .C0(n9), .Y(n49) );
  CLKINVX1 U22 ( .A(n58), .Y(n11) );
  NAND2X1 U23 ( .A(n46), .B(n71), .Y(n38) );
  NAND2X1 U24 ( .A(n30), .B(n5), .Y(n45) );
  NAND2X1 U25 ( .A(n10), .B(n46), .Y(n36) );
  NAND2X1 U26 ( .A(n25), .B(n58), .Y(n33) );
  OAI21XL U27 ( .A0(n15), .A1(n12), .B0(n35), .Y(n48) );
  CLKINVX1 U28 ( .A(n59), .Y(n14) );
  CLKINVX1 U29 ( .A(addr[2]), .Y(n4) );
  OAI31X1 U30 ( .A0(n16), .A1(addr[6]), .A2(n12), .B0(n56), .Y(n55) );
  OAI21XL U31 ( .A0(n30), .A1(n13), .B0(n11), .Y(n56) );
  OAI211X1 U32 ( .A0(n67), .A1(n16), .B0(n45), .C0(n9), .Y(n66) );
  AOI222XL U35 ( .A0(addr[5]), .A1(addr[6]), .B0(n32), .B1(addr[1]), .C0(n6), 
        .C1(n2), .Y(n67) );
  NAND3XL U36 ( .A(n11), .B(n71), .C(addr[4]), .Y(n26) );
  OAI22XL U37 ( .A0(n27), .A1(n28), .B0(n1), .B1(n31), .Y(n65) );
  CLKINVX3 U38 ( .A(addr[4]), .Y(n16) );
  OAI2BB2XL U39 ( .B0(n28), .B1(n37), .A0N(n12), .A1N(n57), .Y(n54) );
  OAI221XL U40 ( .A0(n27), .A1(addr[4]), .B0(n35), .B1(addr[1]), .C0(n26), .Y(
        n57) );
  CLKINVX1 U41 ( .A(addr[6]), .Y(n72) );
  CLKINVX1 U42 ( .A(n62), .Y(n8) );
  OAI21XL U44 ( .A0(n47), .A1(n25), .B0(n50), .Y(n61) );
  NAND3X1 U46 ( .A(n42), .B(n43), .C(n44), .Y(n41) );
  AOI32X1 U47 ( .A0(n47), .A1(n71), .A2(n10), .B0(n11), .B1(n48), .Y(n42) );
  AOI2BB2XL U48 ( .B0(n7), .B1(n22), .A0N(n45), .A1N(addr[5]), .Y(n44) );
  OAI21XL U49 ( .A0(n46), .A1(n13), .B0(n6), .Y(n43) );
  AOI2BB2XL U50 ( .B0(n6), .B1(n20), .A0N(n21), .A1N(n4), .Y(n19) );
  AOI211XL U59 ( .A0(n6), .A1(n22), .B0(n23), .C0(n24), .Y(n21) );
  OAI22XL U60 ( .A0(n27), .A1(n28), .B0(addr[5]), .B1(n29), .Y(n23) );
  CLKINVX1 U61 ( .A(n68), .Y(n9) );
  AOI32XL U62 ( .A0(n10), .A1(n47), .A2(n1), .B0(addr[1]), .B1(n22), .Y(n62)
         );
  AOI222XL U63 ( .A0(n6), .A1(n13), .B0(n22), .B1(n27), .C0(n2), .C1(n70), .Y(
        n63) );
  AOI22XL U64 ( .A0(n65), .A1(n12), .B0(addr[2]), .B1(n66), .Y(n64) );
  NAND2XL U65 ( .A(n32), .B(addr[4]), .Y(n52) );
  AOI211X1 U66 ( .A0(n14), .A1(n33), .B0(n54), .C0(n55), .Y(n53) );
  OAI211X1 U67 ( .A0(n37), .A1(n38), .B0(n39), .C0(n40), .Y(dout[3]) );
  AOI32X1 U68 ( .A0(n2), .A1(n13), .A2(n10), .B0(n49), .B1(n4), .Y(n39) );
  AOI22XL U69 ( .A0(addr[2]), .A1(n41), .B0(n5), .B1(n20), .Y(n40) );
  OAI211X1 U70 ( .A0(addr[2]), .A1(n17), .B0(n18), .C0(n19), .Y(dout[4]) );
  AOI32X1 U71 ( .A0(n11), .A1(n13), .A2(n2), .B0(n3), .B1(n14), .Y(n18) );
  AOI221XL U72 ( .A0(n5), .A1(n32), .B0(n15), .B1(n33), .C0(n34), .Y(n17) );
  CLKINVX3 U73 ( .A(n37), .Y(n6) );
  CLKINVX3 U74 ( .A(addr[1]), .Y(n7) );
  CLKINVX3 U75 ( .A(n47), .Y(n13) );
  CLKINVX3 U76 ( .A(n2), .Y(n71) );
endmodule


module sbox5_0 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n1, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n68, n69, n70;

  OAI222X4 U18 ( .A0(addr[3]), .A1(n32), .B0(n8), .B1(n48), .C0(n13), .C1(n16), 
        .Y(n45) );
  OAI22X2 U40 ( .A0(addr[5]), .A1(n32), .B0(n68), .B1(n24), .Y(n22) );
  NOR2X2 U41 ( .A(n3), .B(addr[3]), .Y(n36) );
  NAND2X2 U45 ( .A(addr[6]), .B(n16), .Y(n24) );
  NAND2X2 U50 ( .A(n16), .B(n8), .Y(n28) );
  NAND2X2 U52 ( .A(addr[1]), .B(n8), .Y(n25) );
  NAND2X2 U54 ( .A(addr[1]), .B(addr[6]), .Y(n32) );
  NAND2X2 U55 ( .A(addr[3]), .B(n13), .Y(n17) );
  CLKINVX1 U1 ( .A(addr[5]), .Y(n1) );
  AOI221XL U2 ( .A0(n45), .A1(n1), .B0(n9), .B1(n14), .C0(n46), .Y(n33) );
  INVX3 U3 ( .A(addr[5]), .Y(n68) );
  OAI221X4 U4 ( .A0(n27), .A1(n28), .B0(n17), .B1(n24), .C0(n29), .Y(n26) );
  OAI221X4 U5 ( .A0(n13), .A1(n24), .B0(n68), .B1(n25), .C0(n18), .Y(n23) );
  OAI221X4 U6 ( .A0(n31), .A1(n17), .B0(n27), .B1(n25), .C0(n53), .Y(n52) );
  OAI31X1 U7 ( .A0(n69), .A1(addr[5]), .A2(addr[1]), .B0(n57), .Y(n65) );
  OAI32X1 U8 ( .A0(n24), .A1(addr[5]), .A2(n3), .B0(n12), .B1(n31), .Y(n59) );
  AOI32XL U9 ( .A0(n14), .A1(n40), .A2(n7), .B0(n2), .B1(n65), .Y(n61) );
  CLKBUFX3 U10 ( .A(addr[4]), .Y(n2) );
  CLKINVX1 U11 ( .A(n57), .Y(n10) );
  NAND2X1 U12 ( .A(n11), .B(n14), .Y(n57) );
  CLKINVX1 U13 ( .A(n28), .Y(n5) );
  CLKXOR2X2 U14 ( .A(n69), .B(n68), .Y(n44) );
  AOI2BB1X1 U15 ( .A0N(n13), .A1N(n1), .B0(n14), .Y(n27) );
  NOR2X1 U16 ( .A(n17), .B(n68), .Y(n47) );
  NOR2BX1 U17 ( .AN(n22), .B(n48), .Y(n55) );
  NAND2X1 U19 ( .A(n5), .B(n68), .Y(n18) );
  CLKINVX1 U20 ( .A(n25), .Y(n7) );
  NAND2X1 U21 ( .A(n7), .B(n68), .Y(n31) );
  CLKINVX1 U22 ( .A(n17), .Y(n12) );
  OAI31X1 U23 ( .A0(n70), .A1(n14), .A2(n25), .B0(n39), .Y(n66) );
  CLKINVX1 U24 ( .A(n32), .Y(n9) );
  OAI2BB2XL U25 ( .B0(n1), .B1(n25), .A0N(n40), .A1N(n11), .Y(n37) );
  CLKINVX1 U26 ( .A(n24), .Y(n11) );
  CLKINVX1 U27 ( .A(n48), .Y(n15) );
  CLKINVX1 U28 ( .A(addr[1]), .Y(n16) );
  CLKINVX1 U29 ( .A(addr[3]), .Y(n69) );
  CLKINVX1 U30 ( .A(addr[6]), .Y(n8) );
  AOI211X1 U31 ( .A0(n47), .A1(addr[1]), .B0(n58), .C0(n59), .Y(n49) );
  OAI2BB2XL U32 ( .B0(n27), .B1(n32), .A0N(n44), .A1N(n5), .Y(n58) );
  AOI211X1 U33 ( .A0(n36), .A1(n54), .B0(n55), .C0(n56), .Y(n53) );
  OAI21XL U34 ( .A0(n8), .A1(n1), .B0(n32), .Y(n54) );
  NOR3XL U35 ( .A(n44), .B(n3), .C(n28), .Y(n56) );
  AOI222XL U36 ( .A0(n9), .A1(n15), .B0(addr[5]), .B1(n30), .C0(n6), .C1(n13), 
        .Y(n29) );
  CLKINVX1 U37 ( .A(n31), .Y(n6) );
  OAI21XL U38 ( .A0(addr[6]), .A1(addr[3]), .B0(n32), .Y(n30) );
  NAND2X1 U39 ( .A(addr[3]), .B(n3), .Y(n48) );
  NAND2X1 U42 ( .A(n2), .B(addr[5]), .Y(n40) );
  NAND2X1 U43 ( .A(n3), .B(n69), .Y(n41) );
  OAI21XL U44 ( .A0(addr[1]), .A1(n41), .B0(n42), .Y(n35) );
  AOI33XL U46 ( .A0(n3), .A1(n43), .A2(addr[5]), .B0(n44), .B1(n13), .B2(
        addr[1]), .Y(n42) );
  OAI21XL U47 ( .A0(n16), .A1(n69), .B0(n24), .Y(n43) );
  OAI21XL U48 ( .A0(addr[6]), .A1(n17), .B0(n39), .Y(n38) );
  NAND2X1 U49 ( .A(n67), .B(n5), .Y(n39) );
  XOR2X1 U51 ( .A(n70), .B(n3), .Y(n67) );
  AOI2BB2XL U53 ( .B0(n36), .B1(n22), .A0N(n2), .A1N(n63), .Y(n62) );
  AOI211X1 U56 ( .A0(n4), .A1(n3), .B0(n64), .C0(n55), .Y(n63) );
  AO22XL U57 ( .A0(n7), .A1(n12), .B0(addr[6]), .B1(n36), .Y(n64) );
  CLKINVX1 U58 ( .A(n18), .Y(n4) );
  CLKINVX1 U59 ( .A(n2), .Y(n70) );
  AO22XL U60 ( .A0(n7), .A1(n15), .B0(addr[6]), .B1(n47), .Y(n46) );
  AOI222XL U61 ( .A0(n22), .A1(n13), .B0(addr[3]), .B1(n23), .C0(n7), .C1(n14), 
        .Y(n21) );
  OAI221X1 U62 ( .A0(n2), .A1(n33), .B0(n28), .B1(n17), .C0(n34), .Y(dout[3])
         );
  AOI222XL U63 ( .A0(n2), .A1(n35), .B0(n36), .B1(n37), .C0(n38), .C1(n1), .Y(
        n34) );
  OAI211X1 U64 ( .A0(n2), .A1(n49), .B0(n50), .C0(n51), .Y(dout[2]) );
  AOI33XL U65 ( .A0(n12), .A1(n40), .A2(n11), .B0(n3), .B1(n44), .B2(n5), .Y(
        n50) );
  AOI222XL U66 ( .A0(n10), .A1(n68), .B0(n2), .B1(n52), .C0(n47), .C1(n9), .Y(
        n51) );
  OAI211X1 U67 ( .A0(n60), .A1(n68), .B0(n61), .C0(n62), .Y(dout[1]) );
  AOI221XL U68 ( .A0(n12), .A1(addr[1]), .B0(n9), .B1(n14), .C0(n66), .Y(n60)
         );
  OAI211X1 U69 ( .A0(n17), .A1(n18), .B0(n19), .C0(n20), .Y(dout[4]) );
  AOI32XL U70 ( .A0(n14), .A1(n24), .A2(addr[5]), .B0(n2), .B1(n26), .Y(n19)
         );
  AOI2BB2X1 U71 ( .B0(n10), .B1(n68), .A0N(n2), .A1N(n21), .Y(n20) );
  BUFX4 U72 ( .A(addr[2]), .Y(n3) );
  CLKINVX3 U73 ( .A(n3), .Y(n13) );
  CLKINVX3 U74 ( .A(n41), .Y(n14) );
endmodule


module sbox6_0 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n81, n82, n83, n84, n85;

  NAND2X2 U39 ( .A(n28), .B(addr[3]), .Y(n19) );
  NOR2X2 U47 ( .A(n83), .B(n81), .Y(n28) );
  NOR2X2 U50 ( .A(n10), .B(n4), .Y(n47) );
  NOR2X2 U58 ( .A(n85), .B(n10), .Y(n41) );
  NAND2X2 U61 ( .A(n69), .B(n63), .Y(n54) );
  NOR2X2 U62 ( .A(n17), .B(addr[1]), .Y(n63) );
  NOR2X2 U63 ( .A(n85), .B(addr[3]), .Y(n69) );
  NAND2X2 U64 ( .A(n49), .B(n35), .Y(n26) );
  NOR2X2 U65 ( .A(n5), .B(addr[3]), .Y(n35) );
  NOR2X2 U66 ( .A(n84), .B(addr[6]), .Y(n49) );
  NOR2X1 U1 ( .A(n83), .B(addr[3]), .Y(n64) );
  AOI211X1 U2 ( .A0(n12), .A1(n10), .B0(n35), .C0(n23), .Y(n45) );
  CLKINVX1 U3 ( .A(n85), .Y(n1) );
  INVX4 U4 ( .A(n4), .Y(n85) );
  CLKBUFX3 U5 ( .A(addr[4]), .Y(n4) );
  CLKINVX1 U6 ( .A(n83), .Y(n2) );
  OAI222X1 U7 ( .A0(n75), .A1(n12), .B0(n5), .B1(n11), .C0(addr[5]), .C1(n8), 
        .Y(n74) );
  BUFX4 U8 ( .A(addr[2]), .Y(n5) );
  OAI221X1 U9 ( .A0(n17), .A1(n9), .B0(n10), .B1(n14), .C0(n80), .Y(n76) );
  INVX2 U10 ( .A(n70), .Y(n14) );
  CLKINVX1 U11 ( .A(addr[3]), .Y(n3) );
  INVX3 U12 ( .A(addr[3]), .Y(n10) );
  OAI221X4 U13 ( .A0(n43), .A1(n16), .B0(n81), .B1(n12), .C0(n13), .Y(n42) );
  NOR2X4 U14 ( .A(addr[1]), .B(addr[6]), .Y(n36) );
  NOR2X4 U15 ( .A(n5), .B(addr[5]), .Y(n23) );
  INVX1 U16 ( .A(n36), .Y(n82) );
  CLKINVX1 U17 ( .A(n41), .Y(n9) );
  NAND2X1 U18 ( .A(n82), .B(n14), .Y(n61) );
  INVXL U19 ( .A(n45), .Y(n6) );
  CLKINVX1 U20 ( .A(n28), .Y(n18) );
  CLKINVX1 U21 ( .A(n49), .Y(n81) );
  CLKINVX1 U22 ( .A(n47), .Y(n8) );
  NOR2X1 U23 ( .A(n14), .B(n43), .Y(n22) );
  NOR2X1 U24 ( .A(n84), .B(n17), .Y(n70) );
  CLKINVX1 U25 ( .A(n63), .Y(n16) );
  OAI211X1 U26 ( .A0(n82), .A1(n9), .B0(n62), .C0(n54), .Y(n58) );
  OAI21XL U27 ( .A0(n63), .A1(n49), .B0(n64), .Y(n62) );
  OAI21XL U28 ( .A0(n34), .A1(n17), .B0(n3), .Y(n80) );
  AOI21X1 U29 ( .A0(n85), .A1(n64), .B0(n41), .Y(n75) );
  OAI2BB2XL U30 ( .B0(n23), .B1(n82), .A0N(n23), .A1N(n49), .Y(n48) );
  CLKINVX1 U31 ( .A(n44), .Y(n13) );
  CLKINVX1 U32 ( .A(n40), .Y(n15) );
  CLKINVX1 U33 ( .A(n69), .Y(n11) );
  NAND2BX1 U34 ( .AN(n22), .B(n29), .Y(n59) );
  CLKINVX1 U35 ( .A(addr[1]), .Y(n84) );
  NOR2X1 U36 ( .A(n14), .B(n2), .Y(n44) );
  NOR2X1 U37 ( .A(addr[1]), .B(n1), .Y(n34) );
  OAI22X1 U38 ( .A0(n8), .A1(n81), .B0(n5), .B1(n15), .Y(n78) );
  NAND2X1 U40 ( .A(n2), .B(n12), .Y(n43) );
  NAND4X1 U41 ( .A(n19), .B(n26), .C(n66), .D(n67), .Y(n65) );
  AOI222XL U42 ( .A0(n68), .A1(n83), .B0(n64), .B1(n36), .C0(n69), .C1(n61), 
        .Y(n67) );
  NAND3X1 U43 ( .A(n5), .B(n8), .C(n70), .Y(n66) );
  OAI221X1 U44 ( .A0(n10), .A1(n16), .B0(n8), .B1(n17), .C0(n15), .Y(n68) );
  AOI22X1 U45 ( .A0(n4), .A1(n51), .B0(addr[5]), .B1(n52), .Y(n37) );
  OAI21XL U46 ( .A0(n45), .A1(n82), .B0(n19), .Y(n51) );
  OAI21XL U48 ( .A0(n53), .A1(n83), .B0(n54), .Y(n52) );
  AOI221XL U49 ( .A0(n47), .A1(n84), .B0(n36), .B1(addr[3]), .C0(n55), .Y(n53)
         );
  OAI22XL U51 ( .A0(n81), .A1(n85), .B0(addr[3]), .B1(n14), .Y(n55) );
  OAI22XL U52 ( .A0(n10), .A1(n17), .B0(addr[1]), .B1(n8), .Y(n24) );
  AOI211X1 U53 ( .A0(n4), .A1(n31), .B0(n32), .C0(n33), .Y(n30) );
  OA21XL U54 ( .A0(n3), .A1(n2), .B0(n34), .Y(n33) );
  OAI2BB2XL U55 ( .B0(n1), .B1(n13), .A0N(n35), .A1N(n36), .Y(n32) );
  OAI22X1 U56 ( .A0(n5), .A1(n81), .B0(n83), .B1(n14), .Y(n31) );
  CLKINVX3 U57 ( .A(addr[5]), .Y(n12) );
  AOI2BB2X1 U59 ( .B0(n5), .B1(n36), .A0N(n2), .A1N(n16), .Y(n29) );
  NOR2X1 U60 ( .A(n16), .B(n1), .Y(n40) );
  AOI2BB2XL U67 ( .B0(n23), .B1(n76), .A0N(n77), .A1N(n12), .Y(n72) );
  AOI211X1 U68 ( .A0(n44), .A1(n4), .B0(n78), .C0(n79), .Y(n77) );
  OAI32X1 U69 ( .A0(n16), .A1(n10), .A2(n83), .B0(n18), .B1(n11), .Y(n79) );
  NAND3X1 U70 ( .A(n19), .B(n26), .C(n27), .Y(n25) );
  AOI32X1 U71 ( .A0(n5), .A1(n84), .A2(n4), .B0(n28), .B1(n85), .Y(n27) );
  AO22XL U72 ( .A0(n23), .A1(n1), .B0(n50), .B1(n85), .Y(n46) );
  OAI21XL U73 ( .A0(n2), .A1(n12), .B0(n43), .Y(n50) );
  CLKINVX1 U74 ( .A(n60), .Y(n7) );
  AOI32XL U75 ( .A0(n61), .A1(n85), .A2(n3), .B0(addr[1]), .B1(n41), .Y(n60)
         );
  OAI211X1 U76 ( .A0(n85), .A1(n26), .B0(n56), .C0(n57), .Y(dout[2]) );
  AOI222XL U77 ( .A0(n58), .A1(n12), .B0(n23), .B1(n7), .C0(n47), .C1(n59), 
        .Y(n57) );
  AOI2BB2XL U78 ( .B0(addr[5]), .B1(n65), .A0N(n83), .A1N(n54), .Y(n56) );
  OAI211X1 U79 ( .A0(n1), .A1(n19), .B0(n20), .C0(n21), .Y(dout[4]) );
  AOI222XL U80 ( .A0(n22), .A1(n10), .B0(n23), .B1(n24), .C0(n25), .C1(n12), 
        .Y(n21) );
  OA22X1 U81 ( .A0(n9), .A1(n29), .B0(n30), .B1(n12), .Y(n20) );
  NAND3X1 U82 ( .A(n37), .B(n38), .C(n39), .Y(dout[3]) );
  AOI32XL U83 ( .A0(n46), .A1(n10), .A2(addr[1]), .B0(n47), .B1(n48), .Y(n38)
         );
  AOI222XL U84 ( .A0(n22), .A1(n85), .B0(n40), .B1(n6), .C0(n41), .C1(n42), 
        .Y(n39) );
  NAND3BX1 U85 ( .AN(n71), .B(n72), .C(n73), .Y(dout[1]) );
  OAI222X1 U86 ( .A0(n26), .A1(n4), .B0(n54), .B1(n83), .C0(n14), .C1(n75), 
        .Y(n71) );
  AOI32XL U87 ( .A0(addr[1]), .A1(n12), .A2(n41), .B0(n36), .B1(n74), .Y(n73)
         );
  CLKINVX3 U88 ( .A(addr[6]), .Y(n17) );
  CLKINVX3 U89 ( .A(n5), .Y(n83) );
endmodule


module sbox7_0 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n83, n84, n85, n86,
         n87;

  OAI222X4 U19 ( .A0(n19), .A1(n41), .B0(n4), .B1(n15), .C0(addr[1]), .C1(n7), 
        .Y(n48) );
  OAI33X4 U33 ( .A0(addr[1]), .A1(n4), .A2(n5), .B0(n16), .B1(n86), .B2(n13), 
        .Y(n73) );
  NOR2X2 U44 ( .A(n87), .B(n4), .Y(n54) );
  NOR2X2 U48 ( .A(addr[1]), .B(addr[6]), .Y(n34) );
  NOR2X2 U51 ( .A(n83), .B(n87), .Y(n45) );
  NOR2X2 U52 ( .A(n16), .B(addr[3]), .Y(n39) );
  NOR2X2 U58 ( .A(n77), .B(n46), .Y(n28) );
  NOR2X2 U60 ( .A(n85), .B(addr[1]), .Y(n77) );
  NOR2X2 U62 ( .A(n11), .B(n3), .Y(n33) );
  NOR2X2 U65 ( .A(n85), .B(n17), .Y(n30) );
  NAND2X1 U1 ( .A(n3), .B(n4), .Y(n51) );
  CLKBUFX3 U2 ( .A(addr[4]), .Y(n4) );
  CLKINVX1 U3 ( .A(n11), .Y(n1) );
  CLKINVX1 U4 ( .A(n86), .Y(n2) );
  CLKBUFX3 U5 ( .A(addr[2]), .Y(n5) );
  OAI22X1 U6 ( .A0(addr[1]), .A1(n7), .B0(n5), .B1(n57), .Y(n70) );
  OAI31X1 U7 ( .A0(n87), .A1(n11), .A2(n17), .B0(n53), .Y(n49) );
  OAI22X1 U8 ( .A0(n4), .A1(n83), .B0(addr[3]), .B1(n10), .Y(n67) );
  NOR2X4 U9 ( .A(n17), .B(addr[6]), .Y(n46) );
  AOI211XL U10 ( .A0(n5), .A1(n14), .B0(n39), .C0(n40), .Y(n38) );
  NOR3XL U11 ( .A(n19), .B(addr[3]), .C(n2), .Y(n40) );
  OAI21XL U12 ( .A0(n3), .A1(n1), .B0(n51), .Y(n81) );
  BUFX4 U13 ( .A(addr[5]), .Y(n3) );
  AOI221XL U14 ( .A0(n30), .A1(n81), .B0(n61), .B1(n14), .C0(n82), .Y(n74) );
  CLKINVX1 U15 ( .A(n30), .Y(n16) );
  OAI2BB2XL U16 ( .B0(n28), .B1(n10), .A0N(n29), .A1N(n30), .Y(n27) );
  CLKINVX1 U17 ( .A(n45), .Y(n21) );
  CLKINVX1 U18 ( .A(n28), .Y(n14) );
  NAND2X1 U20 ( .A(n21), .B(n84), .Y(n65) );
  CLKINVX1 U21 ( .A(n47), .Y(n6) );
  CLKINVX1 U22 ( .A(n61), .Y(n9) );
  NAND2X1 U23 ( .A(n46), .B(n87), .Y(n57) );
  CLKINVX1 U24 ( .A(n33), .Y(n10) );
  NOR2X1 U25 ( .A(n10), .B(n87), .Y(n61) );
  CLKINVX1 U26 ( .A(n34), .Y(n19) );
  OAI22XL U27 ( .A0(n33), .A1(n15), .B0(n17), .B1(n9), .Y(n24) );
  OAI21X1 U28 ( .A0(n11), .A1(n21), .B0(n41), .Y(n29) );
  NAND2X1 U29 ( .A(n54), .B(n83), .Y(n41) );
  CLKINVX1 U30 ( .A(n77), .Y(n18) );
  OAI21XL U31 ( .A0(n51), .A1(n18), .B0(n52), .Y(n50) );
  OAI21XL U32 ( .A0(n45), .A1(n33), .B0(n46), .Y(n52) );
  NOR2X1 U34 ( .A(n83), .B(n7), .Y(n47) );
  CLKINVX1 U35 ( .A(n25), .Y(n7) );
  OAI22XL U36 ( .A0(n33), .A1(n57), .B0(n85), .B1(n6), .Y(n82) );
  CLKINVX1 U37 ( .A(n54), .Y(n13) );
  CLKINVX1 U38 ( .A(n39), .Y(n15) );
  CLKINVX1 U39 ( .A(n36), .Y(n84) );
  NOR2XL U40 ( .A(n45), .B(n11), .Y(n60) );
  CLKINVX1 U41 ( .A(n51), .Y(n12) );
  CLKINVX1 U42 ( .A(n67), .Y(n8) );
  OA21XL U43 ( .A0(n20), .A1(n18), .B0(n53), .Y(n68) );
  CLKINVX1 U45 ( .A(n65), .Y(n20) );
  OAI2BB1XL U46 ( .A0N(n67), .A1N(n46), .B0(n68), .Y(n66) );
  OAI22X1 U47 ( .A0(n83), .A1(n13), .B0(n4), .B1(n84), .Y(n58) );
  NOR4X1 U49 ( .A(n4), .B(addr[3]), .C(n17), .D(n86), .Y(n71) );
  XNOR2X1 U50 ( .A(addr[6]), .B(n5), .Y(n69) );
  AOI211X1 U53 ( .A0(n54), .A1(addr[6]), .B0(n55), .C0(n56), .Y(n42) );
  OAI222X1 U54 ( .A0(n59), .A1(n16), .B0(n60), .B1(n18), .C0(n19), .C1(n9), 
        .Y(n55) );
  OAI2BB2XL U55 ( .B0(n12), .B1(n57), .A0N(n17), .A1N(n58), .Y(n56) );
  OA21XL U56 ( .A0(n87), .A1(n3), .B0(n6), .Y(n59) );
  NAND2X1 U57 ( .A(n5), .B(n34), .Y(n37) );
  CLKINVX1 U59 ( .A(addr[6]), .Y(n85) );
  AOI211X1 U61 ( .A0(n39), .A1(n3), .B0(n78), .C0(n79), .Y(n75) );
  OAI221X1 U63 ( .A0(n17), .A1(n7), .B0(n16), .B1(n10), .C0(n68), .Y(n78) );
  OAI31X1 U64 ( .A0(n87), .A1(n11), .A2(n19), .B0(n80), .Y(n79) );
  AO21XL U66 ( .A0(n51), .A1(n41), .B0(addr[6]), .Y(n80) );
  NOR2X1 U67 ( .A(n11), .B(addr[3]), .Y(n25) );
  AOI21XL U68 ( .A0(addr[3]), .A1(n72), .B0(n73), .Y(n62) );
  OAI2BB1XL U69 ( .A0N(n86), .A1N(n46), .B0(n37), .Y(n72) );
  NAND3X1 U70 ( .A(n34), .B(n87), .C(n3), .Y(n53) );
  NOR2X1 U71 ( .A(addr[3]), .B(n3), .Y(n36) );
  OAI21X1 U72 ( .A0(n5), .A1(n28), .B0(n37), .Y(n32) );
  OAI22XL U73 ( .A0(n28), .A1(n13), .B0(n1), .B1(n38), .Y(n35) );
  AO21X1 U74 ( .A0(n31), .A1(n83), .B0(n32), .Y(n26) );
  OAI21XL U75 ( .A0(n2), .A1(n17), .B0(n18), .Y(n31) );
  OAI221X1 U76 ( .A0(n74), .A1(n86), .B0(n5), .B1(n75), .C0(n76), .Y(dout[1])
         );
  AOI2BB2X1 U77 ( .B0(n77), .B1(n58), .A0N(n37), .A1N(n8), .Y(n76) );
  OAI211X1 U78 ( .A0(n42), .A1(n86), .B0(n43), .C0(n44), .Y(dout[3]) );
  AOI32XL U79 ( .A0(n45), .A1(n1), .A2(n46), .B0(n47), .B1(n34), .Y(n44) );
  OAI31X1 U80 ( .A0(n48), .A1(n49), .A2(n50), .B0(n86), .Y(n43) );
  OAI221X1 U81 ( .A0(n3), .A1(n62), .B0(n63), .B1(n83), .C0(n64), .Y(dout[2])
         );
  AOI32XL U82 ( .A0(n65), .A1(n86), .A2(n30), .B0(n2), .B1(n66), .Y(n64) );
  AOI211X1 U83 ( .A0(n69), .A1(n4), .B0(n70), .C0(n71), .Y(n63) );
  NAND2X1 U84 ( .A(n22), .B(n23), .Y(dout[4]) );
  AOI222XL U85 ( .A0(n34), .A1(n29), .B0(n3), .B1(n35), .C0(n36), .C1(n32), 
        .Y(n22) );
  AOI222XL U86 ( .A0(n5), .A1(n24), .B0(n25), .B1(n26), .C0(n27), .C1(n86), 
        .Y(n23) );
  CLKINVX3 U87 ( .A(n4), .Y(n11) );
  CLKINVX3 U88 ( .A(addr[1]), .Y(n17) );
  CLKINVX3 U89 ( .A(n3), .Y(n83) );
  CLKINVX3 U90 ( .A(n5), .Y(n86) );
  CLKINVX3 U91 ( .A(addr[3]), .Y(n87) );
endmodule


module sbox8_0 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n74, n75;

  NAND2X2 U41 ( .A(addr[6]), .B(n74), .Y(n18) );
  NAND2X2 U48 ( .A(addr[4]), .B(n7), .Y(n26) );
  NAND2X2 U49 ( .A(n2), .B(n4), .Y(n62) );
  NAND2X2 U50 ( .A(addr[1]), .B(n14), .Y(n25) );
  NAND2X2 U54 ( .A(addr[2]), .B(n75), .Y(n33) );
  NAND2X2 U60 ( .A(addr[6]), .B(addr[1]), .Y(n44) );
  NAND2X2 U61 ( .A(n74), .B(n14), .Y(n41) );
  OAI32X1 U1 ( .A0(n14), .A1(addr[4]), .A2(n57), .B0(n34), .B1(n41), .Y(n53)
         );
  OAI31X1 U2 ( .A0(n26), .A1(addr[6]), .A2(n33), .B0(n40), .Y(n39) );
  AOI222X1 U3 ( .A0(n61), .A1(addr[2]), .B0(n4), .B1(n8), .C0(n9), .C1(n57), 
        .Y(n35) );
  OAI222X1 U4 ( .A0(addr[2]), .A1(n23), .B0(n7), .B1(n24), .C0(n25), .C1(n26), 
        .Y(n22) );
  OAI221X1 U5 ( .A0(n44), .A1(n62), .B0(addr[4]), .B1(n41), .C0(n63), .Y(n59)
         );
  NAND2X4 U6 ( .A(addr[4]), .B(n2), .Y(n34) );
  AOI32XL U7 ( .A0(n12), .A1(n10), .A2(n2), .B0(n13), .B1(n32), .Y(n19) );
  OA21XL U8 ( .A0(n9), .A1(n75), .B0(n28), .Y(n71) );
  INVXL U9 ( .A(n30), .Y(n5) );
  INVX3 U10 ( .A(n2), .Y(n7) );
  BUFX4 U11 ( .A(addr[3]), .Y(n2) );
  CLKBUFX3 U12 ( .A(addr[5]), .Y(n1) );
  CLKINVX1 U13 ( .A(n41), .Y(n13) );
  CLKINVX1 U14 ( .A(n42), .Y(n6) );
  CLKINVX1 U15 ( .A(n56), .Y(n3) );
  NAND2X1 U16 ( .A(n7), .B(n4), .Y(n56) );
  NAND2X1 U17 ( .A(n9), .B(n75), .Y(n28) );
  OAI21XL U18 ( .A0(n34), .A1(n75), .B0(n42), .Y(n72) );
  OAI21X1 U19 ( .A0(n4), .A1(n75), .B0(n26), .Y(n61) );
  OAI31XL U20 ( .A0(n34), .A1(n74), .A2(n33), .B0(n31), .Y(n55) );
  CLKINVX1 U21 ( .A(n18), .Y(n16) );
  NAND2X1 U22 ( .A(n10), .B(n7), .Y(n42) );
  OAI22XL U23 ( .A0(n33), .A1(n26), .B0(n10), .B1(n34), .Y(n32) );
  OAI22XL U24 ( .A0(n26), .A1(n41), .B0(n18), .B1(n56), .Y(n54) );
  OAI2BB2XL U25 ( .B0(n34), .B1(n18), .A0N(n61), .A1N(n15), .Y(n60) );
  AOI211XL U26 ( .A0(n41), .A1(n44), .B0(n4), .C0(n28), .Y(n64) );
  CLKINVX1 U27 ( .A(n25), .Y(n12) );
  OAI22XL U28 ( .A0(n10), .A1(n26), .B0(n71), .B1(n62), .Y(n68) );
  NAND2BX2 U29 ( .AN(n71), .B(n7), .Y(n29) );
  NAND2XL U30 ( .A(n34), .B(n56), .Y(n45) );
  OAI2BB2XL U31 ( .B0(n43), .B1(n44), .A0N(n45), .A1N(n12), .Y(n38) );
  NOR2BXL U32 ( .AN(n26), .B(n46), .Y(n43) );
  NAND3X1 U33 ( .A(n45), .B(n74), .C(n10), .Y(n65) );
  AO21X1 U34 ( .A0(n10), .A1(n15), .B0(n48), .Y(n47) );
  OAI33X1 U35 ( .A0(n14), .A1(n7), .A2(n49), .B0(n9), .B1(n46), .B2(n25), .Y(
        n48) );
  OA22XL U36 ( .A0(n42), .A1(n18), .B0(n29), .B1(n25), .Y(n51) );
  CLKINVX1 U37 ( .A(n24), .Y(n11) );
  OAI21XL U38 ( .A0(n12), .A1(n16), .B0(addr[4]), .Y(n63) );
  NAND2X1 U39 ( .A(n1), .B(n9), .Y(n49) );
  OAI221X1 U40 ( .A0(n25), .A1(n28), .B0(addr[1]), .B1(n29), .C0(n5), .Y(n21)
         );
  OAI31XL U42 ( .A0(n9), .A1(n74), .A2(n7), .B0(n31), .Y(n30) );
  NAND2X1 U43 ( .A(n15), .B(addr[2]), .Y(n24) );
  NAND4XL U44 ( .A(n16), .B(n1), .C(n2), .D(addr[2]), .Y(n40) );
  NAND3X1 U45 ( .A(n10), .B(n14), .C(n2), .Y(n31) );
  OAI21XL U46 ( .A0(n1), .A1(n62), .B0(n35), .Y(n73) );
  OAI22XL U47 ( .A0(n41), .A1(n29), .B0(n70), .B1(n49), .Y(n69) );
  AOI221XL U51 ( .A0(n16), .A1(n7), .B0(n15), .B1(n2), .C0(n58), .Y(n70) );
  NOR2X1 U52 ( .A(n1), .B(n2), .Y(n46) );
  NOR2X1 U53 ( .A(n62), .B(addr[6]), .Y(n58) );
  NOR2X1 U55 ( .A(n7), .B(n1), .Y(n57) );
  CLKINVX1 U56 ( .A(n49), .Y(n8) );
  OA21XL U57 ( .A0(n1), .A1(n34), .B0(n29), .Y(n17) );
  AOI221XL U58 ( .A0(n13), .A1(n2), .B0(n15), .B1(addr[4]), .C0(n27), .Y(n23)
         );
  OAI22XL U59 ( .A0(n2), .A1(n74), .B0(addr[4]), .B1(n18), .Y(n27) );
  OAI211X1 U62 ( .A0(addr[2]), .A1(n50), .B0(n51), .C0(n52), .Y(dout[2]) );
  AOI221XL U63 ( .A0(addr[2]), .A1(n53), .B0(n1), .B1(n54), .C0(n55), .Y(n52)
         );
  AOI221XL U64 ( .A0(n58), .A1(n1), .B0(n59), .B1(n75), .C0(n60), .Y(n50) );
  OAI211X1 U65 ( .A0(n17), .A1(n18), .B0(n19), .C0(n20), .Y(dout[4]) );
  AOI222XL U66 ( .A0(n21), .A1(n4), .B0(n1), .B1(n22), .C0(n6), .C1(n15), .Y(
        n20) );
  OAI211X1 U67 ( .A0(addr[1]), .A1(n35), .B0(n36), .C0(n37), .Y(dout[3]) );
  AOI221XL U68 ( .A0(n38), .A1(n9), .B0(n6), .B1(n13), .C0(n39), .Y(n37) );
  AOI2BB2XL U69 ( .B0(n47), .B1(n4), .A0N(n34), .A1N(n24), .Y(n36) );
  NAND4BX1 U70 ( .AN(n64), .B(n65), .C(n66), .D(n67), .Y(dout[1]) );
  AOI221XL U71 ( .A0(n16), .A1(n68), .B0(n3), .B1(n11), .C0(n69), .Y(n67) );
  AOI22X1 U72 ( .A0(n15), .A1(n72), .B0(n12), .B1(n73), .Y(n66) );
  CLKINVX3 U73 ( .A(addr[4]), .Y(n4) );
  CLKINVX3 U74 ( .A(addr[2]), .Y(n9) );
  CLKINVX3 U75 ( .A(n33), .Y(n10) );
  CLKINVX3 U76 ( .A(addr[6]), .Y(n14) );
  CLKINVX3 U77 ( .A(n44), .Y(n15) );
  CLKINVX3 U78 ( .A(addr[1]), .Y(n74) );
  CLKINVX3 U79 ( .A(n1), .Y(n75) );
endmodule


module crp_0 ( P, R, K_sub );
  output [1:32] P;
  input [1:32] R;
  input [1:48] K_sub;
  wire   n1;
  wire   [1:48] X;

  sbox1_0 u0 ( .addr(X[1:6]), .dout({P[9], P[17], P[23], P[31]}) );
  sbox2_0 u1 ( .addr({X[7], n1, X[9:12]}), .dout({P[13], P[28], P[2], P[18]})
         );
  sbox3_0 u2 ( .addr(X[13:18]), .dout({P[24], P[16], P[30], P[6]}) );
  sbox4_0 u3 ( .addr(X[19:24]), .dout({P[26], P[20], P[10], P[1]}) );
  sbox5_0 u4 ( .addr(X[25:30]), .dout({P[8], P[14], P[25], P[3]}) );
  sbox6_0 u5 ( .addr(X[31:36]), .dout({P[4], P[29], P[11], P[19]}) );
  sbox7_0 u6 ( .addr(X[37:42]), .dout({P[32], P[12], P[22], P[7]}) );
  sbox8_0 u7 ( .addr(X[43:48]), .dout({P[5], P[27], P[15], P[21]}) );
  XOR2X1 U1 ( .A(R[1]), .B(K_sub[2]), .Y(X[2]) );
  CLKXOR2X4 U2 ( .A(R[8]), .B(K_sub[11]), .Y(X[11]) );
  CLKXOR2X4 U3 ( .A(R[29]), .B(K_sub[42]), .Y(X[42]) );
  CLKXOR2X4 U4 ( .A(R[5]), .B(K_sub[6]), .Y(X[6]) );
  CLKXOR2X4 U5 ( .A(R[16]), .B(K_sub[25]), .Y(X[25]) );
  CLKXOR2X4 U6 ( .A(R[22]), .B(K_sub[33]), .Y(X[33]) );
  CLKXOR2X4 U7 ( .A(R[29]), .B(K_sub[44]), .Y(X[44]) );
  CLKXOR2X4 U8 ( .A(R[16]), .B(K_sub[23]), .Y(X[23]) );
  CLKXOR2X4 U9 ( .A(R[26]), .B(K_sub[39]), .Y(X[39]) );
  CLKXOR2X4 U10 ( .A(R[10]), .B(K_sub[15]), .Y(X[15]) );
  XNOR2X1 U11 ( .A(R[5]), .B(K_sub[8]), .Y(X[8]) );
  INVX3 U12 ( .A(X[8]), .Y(n1) );
  CLKXOR2X4 U13 ( .A(R[20]), .B(K_sub[31]), .Y(X[31]) );
  CLKXOR2X4 U14 ( .A(R[31]), .B(K_sub[46]), .Y(X[46]) );
  CLKXOR2X4 U15 ( .A(R[12]), .B(K_sub[19]), .Y(X[19]) );
  CLKXOR2X4 U16 ( .A(R[20]), .B(K_sub[29]), .Y(X[29]) );
  CLKXOR2X2 U17 ( .A(R[4]), .B(K_sub[5]), .Y(X[5]) );
  CLKXOR2X2 U18 ( .A(R[15]), .B(K_sub[22]), .Y(X[22]) );
  CLKXOR2X2 U19 ( .A(R[24]), .B(K_sub[35]), .Y(X[35]) );
  CLKXOR2X2 U20 ( .A(R[21]), .B(K_sub[30]), .Y(X[30]) );
  CLKXOR2X2 U21 ( .A(R[12]), .B(K_sub[17]), .Y(X[17]) );
  CLKXOR2X2 U22 ( .A(R[32]), .B(K_sub[1]), .Y(X[1]) );
  CLKXOR2X2 U23 ( .A(R[13]), .B(K_sub[20]), .Y(X[20]) );
  CLKXOR2X2 U24 ( .A(R[18]), .B(K_sub[27]), .Y(X[27]) );
  CLKXOR2X2 U25 ( .A(R[8]), .B(K_sub[13]), .Y(X[13]) );
  CLKXOR2X2 U26 ( .A(R[4]), .B(K_sub[7]), .Y(X[7]) );
  CLKXOR2X2 U27 ( .A(R[24]), .B(K_sub[37]), .Y(X[37]) );
  CLKXOR2X2 U28 ( .A(R[28]), .B(K_sub[43]), .Y(X[43]) );
  CLKXOR2X2 U29 ( .A(R[1]), .B(K_sub[48]), .Y(X[48]) );
  CLKXOR2X2 U30 ( .A(R[17]), .B(K_sub[24]), .Y(X[24]) );
  CLKXOR2X2 U31 ( .A(R[9]), .B(K_sub[12]), .Y(X[12]) );
  CLKXOR2X2 U32 ( .A(R[13]), .B(K_sub[18]), .Y(X[18]) );
  CLKXOR2X2 U33 ( .A(R[25]), .B(K_sub[36]), .Y(X[36]) );
  XOR2X1 U34 ( .A(R[23]), .B(K_sub[34]), .Y(X[34]) );
  XOR2X1 U35 ( .A(R[9]), .B(K_sub[14]), .Y(X[14]) );
  XOR2X1 U36 ( .A(R[30]), .B(K_sub[45]), .Y(X[45]) );
  XOR2X1 U37 ( .A(R[21]), .B(K_sub[32]), .Y(X[32]) );
  XOR2X1 U38 ( .A(R[25]), .B(K_sub[38]), .Y(X[38]) );
  XOR2X1 U39 ( .A(R[27]), .B(K_sub[40]), .Y(X[40]) );
  XOR2X1 U40 ( .A(R[3]), .B(K_sub[4]), .Y(X[4]) );
  XOR2X1 U41 ( .A(R[11]), .B(K_sub[16]), .Y(X[16]) );
  XOR2X1 U42 ( .A(R[7]), .B(K_sub[10]), .Y(X[10]) );
  XOR2X1 U43 ( .A(R[14]), .B(K_sub[21]), .Y(X[21]) );
  XOR2X1 U44 ( .A(R[6]), .B(K_sub[9]), .Y(X[9]) );
  XOR2X1 U45 ( .A(R[2]), .B(K_sub[3]), .Y(X[3]) );
  XOR2X1 U46 ( .A(R[28]), .B(K_sub[41]), .Y(X[41]) );
  XOR2X1 U47 ( .A(R[17]), .B(K_sub[26]), .Y(X[26]) );
  XOR2X1 U48 ( .A(R[32]), .B(K_sub[47]), .Y(X[47]) );
  XOR2X1 U49 ( .A(R[19]), .B(K_sub[28]), .Y(X[28]) );
endmodule


module sbox1_15 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127;

  OAI222X4 U13 ( .A0(addr[5]), .A1(n101), .B0(n1), .B1(n100), .C0(n99), .C1(
        n12), .Y(dout[3]) );
  OAI21X2 U42 ( .A0(n4), .A1(n112), .B0(n106), .Y(n123) );
  NAND2X2 U44 ( .A(addr[6]), .B(n8), .Y(n115) );
  NAND2X2 U48 ( .A(addr[1]), .B(n13), .Y(n114) );
  OAI22X2 U49 ( .A0(n69), .A1(n72), .B0(addr[5]), .B1(n120), .Y(n85) );
  NAND2X2 U50 ( .A(n3), .B(n69), .Y(n120) );
  NOR2X2 U51 ( .A(n69), .B(n3), .Y(n124) );
  NOR2X2 U56 ( .A(n109), .B(n3), .Y(n93) );
  NAND2X2 U57 ( .A(addr[1]), .B(addr[6]), .Y(n109) );
  NAND2X2 U59 ( .A(n8), .B(n13), .Y(n112) );
  NOR2X1 U1 ( .A(n114), .B(n120), .Y(n104) );
  AOI221X4 U2 ( .A0(n7), .A1(n90), .B0(n4), .B1(n93), .C0(n102), .Y(n79) );
  NOR3X1 U3 ( .A(n2), .B(addr[6]), .C(n12), .Y(n102) );
  BUFX4 U4 ( .A(addr[4]), .Y(n2) );
  CLKBUFX3 U5 ( .A(addr[2]), .Y(n1) );
  OAI32X1 U6 ( .A0(n112), .A1(n2), .A2(n4), .B0(n115), .B1(n113), .Y(n80) );
  NOR2BXL U7 ( .AN(n118), .B(n1), .Y(n122) );
  CLKBUFX3 U8 ( .A(addr[2]), .Y(n4) );
  OAI221X4 U9 ( .A0(n88), .A1(n72), .B0(addr[5]), .B1(n87), .C0(n86), .Y(
        dout[2]) );
  OAI221X4 U10 ( .A0(addr[5]), .A1(n127), .B0(n126), .B1(n72), .C0(n125), .Y(
        dout[4]) );
  OA21XL U11 ( .A0(n95), .A1(n115), .B0(n107), .Y(n119) );
  AOI222XL U12 ( .A0(n7), .A1(n1), .B0(n2), .B1(n110), .C0(n9), .C1(n12), .Y(
        n111) );
  AOI2BB2X1 U14 ( .B0(n2), .B1(n9), .A0N(addr[4]), .A1N(n115), .Y(n91) );
  BUFX4 U15 ( .A(addr[3]), .Y(n3) );
  CLKINVX1 U16 ( .A(n112), .Y(n7) );
  CLKINVX1 U17 ( .A(n113), .Y(n11) );
  NAND2BX1 U18 ( .AN(n104), .B(n119), .Y(n84) );
  CLKXOR2X2 U19 ( .A(n70), .B(n12), .Y(n90) );
  NOR2X1 U20 ( .A(n69), .B(n70), .Y(n118) );
  OAI21XL U21 ( .A0(n70), .A1(n114), .B0(n91), .Y(n92) );
  NAND2X1 U22 ( .A(n93), .B(n69), .Y(n107) );
  NAND2X1 U23 ( .A(n12), .B(n70), .Y(n113) );
  OAI211X1 U24 ( .A0(n69), .A1(n114), .B0(n108), .C0(n107), .Y(n89) );
  CLKINVX1 U25 ( .A(n109), .Y(n9) );
  NAND2X1 U26 ( .A(n124), .B(n6), .Y(n108) );
  CLKINVX1 U27 ( .A(n114), .Y(n10) );
  CLKINVX1 U28 ( .A(n115), .Y(n6) );
  CLKINVX1 U29 ( .A(n95), .Y(n71) );
  AO22X1 U30 ( .A0(n90), .A1(n6), .B0(n70), .B1(n123), .Y(n76) );
  OAI31X1 U31 ( .A0(n12), .A1(n3), .A2(n8), .B0(n103), .Y(n105) );
  AOI31XL U32 ( .A0(n8), .A1(n12), .A2(n2), .B0(n102), .Y(n103) );
  CLKINVX1 U33 ( .A(addr[6]), .Y(n13) );
  AOI211X1 U34 ( .A0(n5), .A1(n4), .B0(n117), .C0(n116), .Y(n126) );
  CLKINVX1 U35 ( .A(n108), .Y(n5) );
  AOI211X1 U36 ( .A0(n115), .A1(n114), .B0(n113), .C0(n2), .Y(n116) );
  OAI22X1 U37 ( .A0(n120), .A1(n112), .B0(n111), .B1(n70), .Y(n117) );
  AOI211X1 U38 ( .A0(n9), .A1(n118), .B0(n81), .C0(n80), .Y(n88) );
  OAI22X1 U39 ( .A0(n91), .A1(n12), .B0(n3), .B1(n106), .Y(n81) );
  CLKINVX3 U40 ( .A(addr[5]), .Y(n72) );
  NAND2X1 U41 ( .A(n3), .B(n72), .Y(n95) );
  NAND2X1 U43 ( .A(n10), .B(n1), .Y(n106) );
  XOR2X1 U45 ( .A(n82), .B(n2), .Y(n83) );
  NAND2X1 U46 ( .A(n1), .B(n3), .Y(n82) );
  OAI22XL U47 ( .A0(n3), .A1(n8), .B0(n70), .B1(n112), .Y(n94) );
  AOI211XL U52 ( .A0(n98), .A1(n70), .B0(n97), .C0(n104), .Y(n99) );
  OAI22XL U53 ( .A0(n96), .A1(n69), .B0(n95), .B1(n109), .Y(n97) );
  OAI22XL U54 ( .A0(n13), .A1(n72), .B0(n2), .B1(addr[1]), .Y(n98) );
  AOI221XL U55 ( .A0(n71), .A1(addr[6]), .B0(addr[5]), .B1(n94), .C0(n93), .Y(
        n96) );
  OAI21XL U58 ( .A0(addr[1]), .A1(n120), .B0(n119), .Y(n121) );
  AOI221XL U60 ( .A0(n7), .A1(n118), .B0(n93), .B1(n72), .C0(n75), .Y(n78) );
  OAI31X1 U61 ( .A0(n72), .A1(n2), .A2(n74), .B0(n73), .Y(n75) );
  OA21XL U62 ( .A0(n3), .A1(n13), .B0(n109), .Y(n74) );
  OAI21XL U63 ( .A0(n124), .A1(n85), .B0(n10), .Y(n73) );
  OAI21XL U64 ( .A0(n1), .A1(n8), .B0(n109), .Y(n110) );
  INVX4 U65 ( .A(n4), .Y(n12) );
  AOI222XL U66 ( .A0(n124), .A1(n123), .B0(n122), .B1(addr[6]), .C0(n1), .C1(
        n121), .Y(n125) );
  NOR4BBX1 U67 ( .AN(n107), .BN(n106), .C(n105), .D(n104), .Y(n127) );
  AOI222XL U68 ( .A0(n7), .A1(n90), .B0(n89), .B1(n12), .C0(n123), .C1(n69), 
        .Y(n101) );
  AOI2BB2XL U69 ( .B0(addr[5]), .B1(n92), .A0N(n120), .A1N(addr[1]), .Y(n100)
         );
  AOI32X1 U70 ( .A0(n4), .A1(n85), .A2(n7), .B0(n84), .B1(n12), .Y(n86) );
  AOI222XL U71 ( .A0(n124), .A1(n8), .B0(n83), .B1(addr[1]), .C0(n11), .C1(n13), .Y(n87) );
  OAI221X1 U72 ( .A0(n79), .A1(n72), .B0(n4), .B1(n78), .C0(n77), .Y(dout[1])
         );
  AOI32XL U73 ( .A0(addr[6]), .A1(n85), .A2(n1), .B0(n76), .B1(n72), .Y(n77)
         );
  CLKINVX3 U74 ( .A(addr[1]), .Y(n8) );
  CLKINVX3 U75 ( .A(n2), .Y(n69) );
  CLKINVX3 U76 ( .A(n3), .Y(n70) );
endmodule


module sbox2_15 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147;

  NAND2X2 U55 ( .A(n2), .B(n11), .Y(n136) );
  NAND2X2 U57 ( .A(addr[2]), .B(n9), .Y(n104) );
  NAND2X2 U60 ( .A(addr[5]), .B(addr[2]), .Y(n132) );
  NOR2X2 U61 ( .A(n16), .B(n13), .Y(n101) );
  NAND2X2 U62 ( .A(n15), .B(n82), .Y(n146) );
  NAND2X2 U63 ( .A(n3), .B(n83), .Y(n124) );
  NAND2X2 U64 ( .A(addr[6]), .B(n15), .Y(n122) );
  NAND2X2 U67 ( .A(n3), .B(n2), .Y(n133) );
  AOI222XL U1 ( .A0(n4), .A1(n81), .B0(n88), .B1(n83), .C0(n140), .C1(n13), 
        .Y(n89) );
  CLKINVX1 U2 ( .A(n121), .Y(n16) );
  OAI211X4 U3 ( .A0(n147), .A1(n146), .B0(n145), .C0(n144), .Y(dout[4]) );
  CLKINVX1 U4 ( .A(addr[5]), .Y(n1) );
  INVX3 U5 ( .A(addr[5]), .Y(n9) );
  NAND3XL U6 ( .A(n98), .B(n97), .C(n96), .Y(dout[1]) );
  NAND2X1 U7 ( .A(addr[1]), .B(addr[6]), .Y(n121) );
  CLKINVX2 U8 ( .A(addr[1]), .Y(n15) );
  OAI221X1 U9 ( .A0(addr[1]), .A1(n136), .B0(n133), .B1(n15), .C0(n87), .Y(n95) );
  NOR2X1 U10 ( .A(n104), .B(n2), .Y(n141) );
  NOR2X1 U11 ( .A(n124), .B(n2), .Y(n140) );
  CLKBUFX4 U12 ( .A(addr[4]), .Y(n2) );
  NAND2X4 U13 ( .A(addr[1]), .B(n82), .Y(n114) );
  INVX3 U14 ( .A(addr[6]), .Y(n82) );
  NAND2XL U15 ( .A(n102), .B(n11), .Y(n109) );
  AOI211XL U16 ( .A0(n10), .A1(n95), .B0(n94), .C0(n93), .Y(n96) );
  AOI2BB2X1 U17 ( .B0(n9), .B1(n12), .A0N(n104), .A1N(n136), .Y(n117) );
  NOR3BXL U18 ( .AN(n135), .B(n134), .C(n4), .Y(n147) );
  BUFX4 U19 ( .A(addr[3]), .Y(n3) );
  NAND2X1 U20 ( .A(n4), .B(n16), .Y(n113) );
  CLKINVX1 U21 ( .A(n146), .Y(n13) );
  CLKINVX1 U22 ( .A(n115), .Y(n4) );
  CLKINVX1 U23 ( .A(n122), .Y(n14) );
  OAI31X1 U24 ( .A0(n124), .A1(n82), .A2(n9), .B0(n123), .Y(n128) );
  OAI21XL U25 ( .A0(n9), .A1(n15), .B0(n140), .Y(n123) );
  OAI22X1 U26 ( .A0(n122), .A1(n124), .B0(n101), .B1(n132), .Y(n84) );
  INVX1 U27 ( .A(n114), .Y(n81) );
  OAI22X1 U28 ( .A0(n122), .A1(n11), .B0(n5), .B1(n121), .Y(n129) );
  NAND3X1 U29 ( .A(n5), .B(n9), .C(n15), .Y(n111) );
  NAND2X1 U30 ( .A(n11), .B(n5), .Y(n115) );
  OAI21XL U31 ( .A0(n83), .A1(n133), .B0(n135), .Y(n85) );
  OAI22XL U32 ( .A0(n117), .A1(n146), .B0(n116), .B1(n132), .Y(n118) );
  AOI222XL U33 ( .A0(n81), .A1(n115), .B0(n6), .B1(n82), .C0(n4), .C1(n13), 
        .Y(n116) );
  CLKINVX1 U34 ( .A(n104), .Y(n8) );
  OAI2BB2XL U35 ( .B0(n114), .B1(n135), .A0N(n126), .A1N(n6), .Y(n106) );
  OAI21XL U36 ( .A0(n112), .A1(n114), .B0(n111), .Y(n120) );
  OAI21XL U37 ( .A0(n133), .A1(n114), .B0(n113), .Y(n119) );
  CLKINVX1 U38 ( .A(n124), .Y(n12) );
  CLKINVX1 U39 ( .A(n136), .Y(n7) );
  CLKINVX1 U40 ( .A(n133), .Y(n6) );
  CLKINVX1 U41 ( .A(n132), .Y(n10) );
  AOI2BB1X1 U42 ( .A0N(n126), .A1N(n125), .B0(n136), .Y(n127) );
  OAI22XL U43 ( .A0(n104), .A1(n114), .B0(n101), .B1(n132), .Y(n102) );
  AO21XL U44 ( .A0(n83), .A1(n7), .B0(n141), .Y(n86) );
  AO21X1 U45 ( .A0(n11), .A1(n8), .B0(n140), .Y(n142) );
  NAND3X1 U46 ( .A(n83), .B(n5), .C(addr[5]), .Y(n135) );
  OAI22X1 U47 ( .A0(addr[5]), .A1(n121), .B0(n122), .B1(n9), .Y(n126) );
  AOI2BB1X1 U48 ( .A0N(n3), .A1N(n1), .B0(n7), .Y(n112) );
  NOR3X1 U49 ( .A(addr[1]), .B(addr[2]), .C(n9), .Y(n125) );
  AOI2BB1XL U50 ( .A0N(n92), .A1N(n91), .B0(addr[5]), .Y(n93) );
  OAI22XL U51 ( .A0(n117), .A1(n114), .B0(n89), .B1(n1), .Y(n94) );
  OAI31XL U52 ( .A0(n114), .A1(n2), .A2(n11), .B0(n90), .Y(n91) );
  OAI21XL U53 ( .A0(n6), .A1(n12), .B0(n14), .Y(n90) );
  NAND2X1 U54 ( .A(n81), .B(n2), .Y(n137) );
  OAI31XL U56 ( .A0(n101), .A1(n3), .A2(addr[2]), .B0(n113), .Y(n92) );
  OAI211X1 U58 ( .A0(n139), .A1(n9), .B0(n138), .C0(n137), .Y(n143) );
  NAND3X1 U59 ( .A(n5), .B(n9), .C(addr[6]), .Y(n138) );
  AOI2BB2X1 U65 ( .B0(n14), .B1(n11), .A0N(n15), .A1N(n136), .Y(n139) );
  OAI22XL U66 ( .A0(addr[5]), .A1(n133), .B0(n3), .B1(n132), .Y(n134) );
  OAI2BB2XL U68 ( .B0(n112), .B1(n122), .A0N(n1), .A1N(n99), .Y(n100) );
  OAI211X1 U69 ( .A0(n146), .A1(n2), .B0(n137), .C0(n113), .Y(n99) );
  NAND3X1 U70 ( .A(n14), .B(n5), .C(n3), .Y(n87) );
  AOI2BB2XL U71 ( .B0(n3), .B1(n105), .A0N(n137), .A1N(n132), .Y(n108) );
  OAI211XL U72 ( .A0(n104), .A1(n146), .B0(n103), .C0(n111), .Y(n105) );
  NAND3XL U73 ( .A(addr[5]), .B(n5), .C(n16), .Y(n103) );
  OAI22XL U74 ( .A0(n3), .A1(n114), .B0(n82), .B1(n115), .Y(n88) );
  NAND4X1 U75 ( .A(n110), .B(n109), .C(n108), .D(n107), .Y(dout[2]) );
  AOI32XL U76 ( .A0(addr[1]), .A1(addr[2]), .A2(n7), .B0(n100), .B1(n83), .Y(
        n110) );
  AOI221XL U77 ( .A0(n125), .A1(addr[4]), .B0(n141), .B1(n14), .C0(n106), .Y(
        n107) );
  AOI33XL U78 ( .A0(n14), .A1(n8), .A2(n2), .B0(n10), .B1(n146), .B2(n3), .Y(
        n145) );
  AOI222XL U79 ( .A0(n143), .A1(n83), .B0(n16), .B1(n142), .C0(n81), .C1(n141), 
        .Y(n144) );
  AOI32XL U80 ( .A0(n8), .A1(n15), .A2(n4), .B0(n13), .B1(n86), .Y(n97) );
  AOI22X1 U81 ( .A0(n16), .A1(n85), .B0(n2), .B1(n84), .Y(n98) );
  NAND2X1 U82 ( .A(n131), .B(n130), .Y(dout[3]) );
  AOI221XL U83 ( .A0(n120), .A1(n83), .B0(addr[2]), .B1(n119), .C0(n118), .Y(
        n131) );
  AOI211X1 U84 ( .A0(n8), .A1(n129), .B0(n128), .C0(n127), .Y(n130) );
  CLKINVX3 U85 ( .A(n2), .Y(n5) );
  CLKINVX3 U86 ( .A(n3), .Y(n11) );
  CLKINVX3 U87 ( .A(addr[2]), .Y(n83) );
endmodule


module sbox3_15 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133;

  NOR2X2 U35 ( .A(n15), .B(addr[3]), .Y(n108) );
  NOR2X2 U50 ( .A(addr[1]), .B(addr[6]), .Y(n107) );
  NOR2X2 U52 ( .A(n20), .B(n2), .Y(n87) );
  NOR2X2 U56 ( .A(n20), .B(n77), .Y(n94) );
  NOR2X1 U1 ( .A(n15), .B(n20), .Y(n106) );
  OAI221X1 U2 ( .A0(n124), .A1(n15), .B0(n3), .B1(addr[1]), .C0(n13), .Y(n104)
         );
  OAI22XL U3 ( .A0(n2), .A1(n77), .B0(n3), .B1(n14), .Y(n123) );
  BUFX4 U4 ( .A(addr[4]), .Y(n2) );
  CLKBUFX3 U5 ( .A(n77), .Y(n1) );
  OAI33X1 U6 ( .A0(n17), .A1(n125), .A2(n77), .B0(n15), .B1(n94), .B2(n119), 
        .Y(n79) );
  INVX3 U7 ( .A(n3), .Y(n77) );
  NOR2X1 U8 ( .A(n9), .B(n3), .Y(n91) );
  NOR2X1 U9 ( .A(n17), .B(n3), .Y(n121) );
  NOR2X1 U10 ( .A(n13), .B(n3), .Y(n95) );
  NOR2X1 U11 ( .A(n3), .B(n2), .Y(n110) );
  CLKBUFX4 U12 ( .A(addr[2]), .Y(n3) );
  OAI221X1 U13 ( .A0(addr[5]), .A1(n90), .B0(n89), .B1(n78), .C0(n88), .Y(
        dout[1]) );
  NOR2X4 U14 ( .A(n10), .B(n76), .Y(n124) );
  NOR2X4 U15 ( .A(addr[3]), .B(n2), .Y(n130) );
  NOR2X4 U16 ( .A(n76), .B(addr[6]), .Y(n125) );
  INVX3 U17 ( .A(addr[1]), .Y(n76) );
  NAND2XL U18 ( .A(n94), .B(n124), .Y(n132) );
  OAI211XL U19 ( .A0(n2), .A1(n8), .B0(n128), .C0(n127), .Y(n129) );
  NAND4XL U20 ( .A(n114), .B(n113), .C(n112), .D(n111), .Y(n115) );
  CLKINVX1 U21 ( .A(n132), .Y(n6) );
  INVX1 U22 ( .A(n124), .Y(n4) );
  CLKINVX1 U23 ( .A(n106), .Y(n14) );
  NAND2X1 U24 ( .A(n9), .B(n11), .Y(n122) );
  CLKINVX1 U25 ( .A(n86), .Y(n11) );
  CLKINVX1 U26 ( .A(n120), .Y(n19) );
  CLKINVX1 U27 ( .A(n119), .Y(n5) );
  CLKINVX1 U28 ( .A(n114), .Y(n7) );
  CLKINVX1 U29 ( .A(n107), .Y(n13) );
  NOR2X1 U30 ( .A(n9), .B(n77), .Y(n103) );
  NOR2X1 U31 ( .A(n4), .B(n77), .Y(n109) );
  INVX1 U32 ( .A(n125), .Y(n12) );
  AOI21X1 U33 ( .A0(n20), .A1(n77), .B0(n94), .Y(n120) );
  OAI21XL U34 ( .A0(n110), .A1(n130), .B0(n124), .Y(n82) );
  CLKINVX1 U36 ( .A(n81), .Y(n9) );
  NOR2X1 U37 ( .A(n12), .B(n15), .Y(n86) );
  NOR2X1 U38 ( .A(n124), .B(n107), .Y(n119) );
  OAI21XL U39 ( .A0(n109), .A1(n91), .B0(n130), .Y(n100) );
  NAND2X1 U40 ( .A(n103), .B(n87), .Y(n114) );
  CLKINVX1 U41 ( .A(n87), .Y(n17) );
  CLKINVX1 U42 ( .A(n91), .Y(n8) );
  CLKINVX1 U43 ( .A(n110), .Y(n18) );
  CLKINVX1 U44 ( .A(n121), .Y(n16) );
  OR2X1 U45 ( .A(n103), .B(n95), .Y(n126) );
  OAI221X1 U46 ( .A0(n12), .A1(n18), .B0(n77), .B1(n11), .C0(n93), .Y(n98) );
  AOI221XL U47 ( .A0(n95), .A1(n2), .B0(n92), .B1(n15), .C0(n6), .Y(n93) );
  OAI21XL U48 ( .A0(n1), .A1(n13), .B0(n8), .Y(n92) );
  XNOR2X1 U49 ( .A(addr[5]), .B(addr[3]), .Y(n102) );
  CLKINVX1 U51 ( .A(addr[5]), .Y(n78) );
  OAI221X1 U53 ( .A0(n13), .A1(n18), .B0(n4), .B1(n17), .C0(n105), .Y(n116) );
  AOI221XL U54 ( .A0(addr[3]), .A1(n104), .B0(n103), .B1(n130), .C0(n6), .Y(
        n105) );
  CLKINVX1 U55 ( .A(addr[6]), .Y(n10) );
  NAND3X1 U57 ( .A(n3), .B(n76), .C(n108), .Y(n113) );
  NOR2X1 U58 ( .A(n10), .B(addr[1]), .Y(n81) );
  AOI32XL U59 ( .A0(n1), .A1(n20), .A2(n124), .B0(n123), .B1(n10), .Y(n128) );
  AOI22XL U60 ( .A0(n2), .A1(n126), .B0(n125), .B1(n130), .Y(n127) );
  AOI222XL U61 ( .A0(n110), .A1(n125), .B0(n109), .B1(n20), .C0(n108), .C1(
        n107), .Y(n111) );
  OAI211XL U62 ( .A0(n106), .A1(n130), .B0(n1), .C0(addr[6]), .Y(n112) );
  OAI21XL U63 ( .A0(n3), .A1(addr[1]), .B0(n12), .Y(n80) );
  AOI221XL U64 ( .A0(n86), .A1(n20), .B0(n87), .B1(n125), .C0(n85), .Y(n89) );
  OAI211X1 U65 ( .A0(n84), .A1(n77), .B0(n83), .C0(n82), .Y(n85) );
  AOI222XL U66 ( .A0(n81), .A1(n20), .B0(n107), .B1(n106), .C0(n130), .C1(n76), 
        .Y(n84) );
  OAI21XL U67 ( .A0(n91), .A1(n6), .B0(addr[4]), .Y(n83) );
  AOI221XL U68 ( .A0(n125), .A1(n19), .B0(addr[3]), .B1(n126), .C0(n96), .Y(
        n97) );
  OAI22X1 U69 ( .A0(n4), .A1(n16), .B0(n14), .B1(n9), .Y(n96) );
  OAI211X1 U70 ( .A0(n13), .A1(n16), .B0(n118), .C0(n117), .Y(dout[3]) );
  AOI32XL U71 ( .A0(n125), .A1(n3), .A2(n102), .B0(n108), .B1(n109), .Y(n118)
         );
  AOI22XL U72 ( .A0(n116), .A1(n78), .B0(addr[5]), .B1(n115), .Y(n117) );
  AOI221XL U73 ( .A0(n121), .A1(n125), .B0(n95), .B1(n108), .C0(n7), .Y(n88)
         );
  AOI221XL U74 ( .A0(n130), .A1(n80), .B0(n94), .B1(n122), .C0(n79), .Y(n90)
         );
  NAND4X1 U75 ( .A(n101), .B(n113), .C(n100), .D(n99), .Y(dout[2]) );
  NAND3XL U76 ( .A(n2), .B(n124), .C(n102), .Y(n101) );
  AOI2BB2XL U77 ( .B0(addr[5]), .B1(n98), .A0N(addr[5]), .A1N(n97), .Y(n99) );
  OAI221X1 U78 ( .A0(n133), .A1(n78), .B0(n2), .B1(n132), .C0(n131), .Y(
        dout[4]) );
  AOI32XL U79 ( .A0(n130), .A1(n10), .A2(addr[2]), .B0(n129), .B1(n78), .Y(
        n131) );
  AOI222XL U80 ( .A0(n19), .A1(n122), .B0(n121), .B1(addr[1]), .C0(n120), .C1(
        n5), .Y(n133) );
  CLKINVX3 U81 ( .A(n2), .Y(n15) );
  CLKINVX3 U82 ( .A(addr[3]), .Y(n20) );
endmodule


module sbox4_15 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126;

  OAI32X4 U12 ( .A0(n12), .A1(n2), .A2(addr[2]), .B0(n11), .B1(n108), .Y(n123)
         );
  OAI222X4 U20 ( .A0(addr[2]), .A1(n92), .B0(n106), .B1(n91), .C0(n90), .C1(
        n14), .Y(dout[2]) );
  OAI222X4 U33 ( .A0(addr[4]), .A1(n106), .B0(n6), .B1(n108), .C0(n2), .C1(
        n118), .Y(n83) );
  NAND2X2 U34 ( .A(addr[4]), .B(n2), .Y(n108) );
  NOR2X2 U43 ( .A(n72), .B(addr[4]), .Y(n113) );
  NOR2X2 U45 ( .A(n11), .B(n2), .Y(n111) );
  NAND2X2 U51 ( .A(n6), .B(n71), .Y(n118) );
  NOR2X2 U52 ( .A(n16), .B(addr[5]), .Y(n97) );
  NAND2X2 U53 ( .A(addr[6]), .B(addr[1]), .Y(n85) );
  NAND2X2 U54 ( .A(addr[1]), .B(n71), .Y(n116) );
  NOR2X2 U55 ( .A(n115), .B(n11), .Y(n121) );
  NAND2X2 U56 ( .A(n72), .B(n16), .Y(n115) );
  NAND2X2 U57 ( .A(addr[5]), .B(n16), .Y(n96) );
  NAND2X2 U58 ( .A(addr[6]), .B(n6), .Y(n106) );
  OAI222X1 U1 ( .A0(n12), .A1(n85), .B0(n97), .B1(n116), .C0(n16), .C1(n118), 
        .Y(n73) );
  CLKINVX1 U2 ( .A(n116), .Y(n9) );
  OAI31X4 U3 ( .A0(n118), .A1(n11), .A2(n16), .B0(n117), .Y(n119) );
  CLKINVX1 U4 ( .A(n72), .Y(n1) );
  CLKBUFX3 U5 ( .A(addr[3]), .Y(n2) );
  OAI221X1 U6 ( .A0(addr[2]), .A1(n80), .B0(n118), .B1(n105), .C0(n79), .Y(
        dout[1]) );
  INVX4 U7 ( .A(addr[5]), .Y(n11) );
  OAI31X1 U8 ( .A0(n108), .A1(addr[5]), .A2(n5), .B0(n107), .Y(n109) );
  AOI222XL U9 ( .A0(n16), .A1(n71), .B0(n113), .B1(n6), .C0(addr[1]), .C1(n72), 
        .Y(n114) );
  OAI222X1 U10 ( .A0(addr[1]), .A1(n84), .B0(n85), .B1(n74), .C0(n72), .C1(
        n107), .Y(n75) );
  NAND2XL U11 ( .A(n1), .B(addr[5]), .Y(n84) );
  AOI211XL U13 ( .A0(n83), .A1(n11), .B0(n82), .C0(n7), .Y(n92) );
  NAND2XL U14 ( .A(n16), .B(n11), .Y(n74) );
  CLKINVX1 U15 ( .A(n118), .Y(n3) );
  CLKINVX1 U16 ( .A(n115), .Y(n15) );
  CLKINVX1 U17 ( .A(n112), .Y(n4) );
  OAI21X1 U18 ( .A0(n9), .A1(n5), .B0(n14), .Y(n112) );
  AOI22X1 U19 ( .A0(n10), .A1(n111), .B0(n5), .B1(n113), .Y(n93) );
  OAI211X1 U21 ( .A0(n6), .A1(n115), .B0(n93), .C0(n8), .Y(n94) );
  CLKINVX1 U22 ( .A(n85), .Y(n10) );
  NAND2X1 U23 ( .A(n97), .B(n72), .Y(n105) );
  NAND2X1 U24 ( .A(n113), .B(n3), .Y(n98) );
  NAND2X1 U25 ( .A(n9), .B(n97), .Y(n107) );
  NAND2X1 U26 ( .A(n118), .B(n85), .Y(n110) );
  OAI21XL U27 ( .A0(n15), .A1(n11), .B0(n108), .Y(n95) );
  CLKINVX1 U28 ( .A(n84), .Y(n13) );
  CLKINVX1 U29 ( .A(addr[2]), .Y(n14) );
  OAI31X1 U30 ( .A0(n16), .A1(addr[6]), .A2(n11), .B0(n87), .Y(n88) );
  OAI21XL U31 ( .A0(n113), .A1(n12), .B0(n10), .Y(n87) );
  OAI211X1 U32 ( .A0(n76), .A1(n16), .B0(n98), .C0(n8), .Y(n77) );
  AOI222XL U35 ( .A0(addr[5]), .A1(addr[6]), .B0(n111), .B1(addr[1]), .C0(n5), 
        .C1(n2), .Y(n76) );
  NAND3XL U36 ( .A(n10), .B(n72), .C(addr[4]), .Y(n117) );
  OAI22XL U37 ( .A0(n116), .A1(n115), .B0(n1), .B1(n112), .Y(n78) );
  CLKINVX3 U38 ( .A(addr[4]), .Y(n16) );
  OAI2BB2XL U39 ( .B0(n115), .B1(n106), .A0N(n11), .A1N(n86), .Y(n89) );
  OAI221XL U40 ( .A0(n116), .A1(addr[4]), .B0(n108), .B1(addr[1]), .C0(n117), 
        .Y(n86) );
  CLKINVX1 U41 ( .A(addr[6]), .Y(n71) );
  CLKINVX1 U42 ( .A(n81), .Y(n7) );
  OAI21XL U44 ( .A0(n96), .A1(n118), .B0(n93), .Y(n82) );
  NAND3X1 U46 ( .A(n101), .B(n100), .C(n99), .Y(n102) );
  AOI32X1 U47 ( .A0(n96), .A1(n72), .A2(n9), .B0(n10), .B1(n95), .Y(n101) );
  AOI2BB2XL U48 ( .B0(n6), .B1(n121), .A0N(n98), .A1N(addr[5]), .Y(n99) );
  OAI21XL U49 ( .A0(n97), .A1(n12), .B0(n5), .Y(n100) );
  AOI2BB2XL U50 ( .B0(n5), .B1(n123), .A0N(n122), .A1N(n14), .Y(n124) );
  AOI211XL U59 ( .A0(n5), .A1(n121), .B0(n120), .C0(n119), .Y(n122) );
  OAI22XL U60 ( .A0(n116), .A1(n115), .B0(addr[5]), .B1(n114), .Y(n120) );
  CLKINVX1 U61 ( .A(n75), .Y(n8) );
  AOI32XL U62 ( .A0(n9), .A1(n96), .A2(n1), .B0(addr[1]), .B1(n121), .Y(n81)
         );
  AOI222XL U63 ( .A0(n5), .A1(n12), .B0(n121), .B1(n116), .C0(n2), .C1(n73), 
        .Y(n80) );
  AOI22XL U64 ( .A0(n78), .A1(n11), .B0(addr[2]), .B1(n77), .Y(n79) );
  NAND2XL U65 ( .A(n111), .B(addr[4]), .Y(n91) );
  AOI211X1 U66 ( .A0(n13), .A1(n110), .B0(n89), .C0(n88), .Y(n90) );
  OAI211X1 U67 ( .A0(n106), .A1(n105), .B0(n104), .C0(n103), .Y(dout[3]) );
  AOI32X1 U68 ( .A0(n2), .A1(n12), .A2(n9), .B0(n94), .B1(n14), .Y(n104) );
  AOI22XL U69 ( .A0(addr[2]), .A1(n102), .B0(n3), .B1(n123), .Y(n103) );
  OAI211X1 U70 ( .A0(addr[2]), .A1(n126), .B0(n125), .C0(n124), .Y(dout[4]) );
  AOI32X1 U71 ( .A0(n10), .A1(n12), .A2(n2), .B0(n4), .B1(n13), .Y(n125) );
  AOI221XL U72 ( .A0(n3), .A1(n111), .B0(n15), .B1(n110), .C0(n109), .Y(n126)
         );
  CLKINVX3 U73 ( .A(n106), .Y(n5) );
  CLKINVX3 U74 ( .A(addr[1]), .Y(n6) );
  CLKINVX3 U75 ( .A(n96), .Y(n12) );
  CLKINVX3 U76 ( .A(n2), .Y(n72) );
endmodule


module sbox5_15 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121;

  OAI222X4 U18 ( .A0(addr[3]), .A1(n106), .B0(n68), .B1(n90), .C0(n6), .C1(n13), .Y(n93) );
  OAI22X2 U40 ( .A0(addr[5]), .A1(n106), .B0(n69), .B1(n114), .Y(n116) );
  NOR2X2 U41 ( .A(n3), .B(addr[3]), .Y(n102) );
  NAND2X2 U45 ( .A(addr[6]), .B(n13), .Y(n114) );
  NAND2X2 U50 ( .A(n13), .B(n68), .Y(n110) );
  NAND2X2 U52 ( .A(addr[1]), .B(n68), .Y(n113) );
  NAND2X2 U54 ( .A(addr[1]), .B(addr[6]), .Y(n106) );
  NAND2X2 U55 ( .A(addr[3]), .B(n6), .Y(n121) );
  OAI221X4 U1 ( .A0(n111), .A1(n110), .B0(n121), .B1(n114), .C0(n109), .Y(n112) );
  OAI221X4 U2 ( .A0(n107), .A1(n121), .B0(n111), .B1(n113), .C0(n85), .Y(n86)
         );
  OAI31X1 U3 ( .A0(n70), .A1(addr[5]), .A2(addr[1]), .B0(n81), .Y(n73) );
  CLKINVX1 U4 ( .A(addr[5]), .Y(n1) );
  OAI221X4 U5 ( .A0(n6), .A1(n114), .B0(n69), .B1(n113), .C0(n120), .Y(n115)
         );
  AOI221XL U6 ( .A0(n93), .A1(n1), .B0(n14), .B1(n8), .C0(n92), .Y(n105) );
  INVX3 U7 ( .A(addr[5]), .Y(n69) );
  OAI32X1 U8 ( .A0(n114), .A1(addr[5]), .A2(n3), .B0(n5), .B1(n107), .Y(n79)
         );
  AOI32XL U9 ( .A0(n8), .A1(n98), .A2(n16), .B0(n2), .B1(n73), .Y(n77) );
  CLKBUFX3 U10 ( .A(addr[4]), .Y(n2) );
  CLKINVX1 U11 ( .A(n81), .Y(n7) );
  NAND2X1 U12 ( .A(n10), .B(n8), .Y(n81) );
  CLKINVX1 U13 ( .A(n110), .Y(n12) );
  CLKXOR2X2 U14 ( .A(n70), .B(n69), .Y(n94) );
  AOI2BB1X1 U15 ( .A0N(n6), .A1N(n1), .B0(n8), .Y(n111) );
  NOR2X1 U16 ( .A(n121), .B(n69), .Y(n91) );
  NOR2BX1 U17 ( .AN(n116), .B(n90), .Y(n83) );
  NAND2X1 U19 ( .A(n12), .B(n69), .Y(n120) );
  CLKINVX1 U20 ( .A(n113), .Y(n16) );
  NAND2X1 U21 ( .A(n16), .B(n69), .Y(n107) );
  CLKINVX1 U22 ( .A(n121), .Y(n5) );
  OAI31X1 U23 ( .A0(n4), .A1(n8), .A2(n113), .B0(n99), .Y(n72) );
  CLKINVX1 U24 ( .A(n106), .Y(n14) );
  OAI2BB2XL U25 ( .B0(n1), .B1(n113), .A0N(n98), .A1N(n10), .Y(n101) );
  CLKINVX1 U26 ( .A(n114), .Y(n10) );
  CLKINVX1 U27 ( .A(n90), .Y(n9) );
  CLKINVX1 U28 ( .A(addr[1]), .Y(n13) );
  CLKINVX1 U29 ( .A(addr[3]), .Y(n70) );
  CLKINVX1 U30 ( .A(addr[6]), .Y(n68) );
  AOI211X1 U31 ( .A0(n91), .A1(addr[1]), .B0(n80), .C0(n79), .Y(n89) );
  OAI2BB2XL U32 ( .B0(n111), .B1(n106), .A0N(n94), .A1N(n12), .Y(n80) );
  AOI211X1 U33 ( .A0(n102), .A1(n84), .B0(n83), .C0(n82), .Y(n85) );
  OAI21XL U34 ( .A0(n68), .A1(n1), .B0(n106), .Y(n84) );
  NOR3XL U35 ( .A(n94), .B(n3), .C(n110), .Y(n82) );
  AOI222XL U36 ( .A0(n14), .A1(n9), .B0(addr[5]), .B1(n108), .C0(n15), .C1(n6), 
        .Y(n109) );
  CLKINVX1 U37 ( .A(n107), .Y(n15) );
  OAI21XL U38 ( .A0(addr[6]), .A1(addr[3]), .B0(n106), .Y(n108) );
  NAND2X1 U39 ( .A(addr[3]), .B(n3), .Y(n90) );
  NAND2X1 U42 ( .A(n2), .B(addr[5]), .Y(n98) );
  NAND2X1 U43 ( .A(n3), .B(n70), .Y(n97) );
  OAI21XL U44 ( .A0(addr[1]), .A1(n97), .B0(n96), .Y(n103) );
  AOI33XL U46 ( .A0(n3), .A1(n95), .A2(addr[5]), .B0(n94), .B1(n6), .B2(
        addr[1]), .Y(n96) );
  OAI21XL U47 ( .A0(n13), .A1(n70), .B0(n114), .Y(n95) );
  OAI21XL U48 ( .A0(addr[6]), .A1(n121), .B0(n99), .Y(n100) );
  NAND2X1 U49 ( .A(n71), .B(n12), .Y(n99) );
  XOR2X1 U51 ( .A(n4), .B(n3), .Y(n71) );
  AOI2BB2XL U53 ( .B0(n102), .B1(n116), .A0N(n2), .A1N(n75), .Y(n76) );
  AOI211X1 U56 ( .A0(n11), .A1(n3), .B0(n74), .C0(n83), .Y(n75) );
  AO22XL U57 ( .A0(n16), .A1(n5), .B0(addr[6]), .B1(n102), .Y(n74) );
  CLKINVX1 U58 ( .A(n120), .Y(n11) );
  CLKINVX1 U59 ( .A(n2), .Y(n4) );
  AO22XL U60 ( .A0(n16), .A1(n9), .B0(addr[6]), .B1(n91), .Y(n92) );
  AOI222XL U61 ( .A0(n116), .A1(n6), .B0(addr[3]), .B1(n115), .C0(n16), .C1(n8), .Y(n117) );
  OAI221X1 U62 ( .A0(n2), .A1(n105), .B0(n110), .B1(n121), .C0(n104), .Y(
        dout[3]) );
  AOI222XL U63 ( .A0(n2), .A1(n103), .B0(n102), .B1(n101), .C0(n100), .C1(n1), 
        .Y(n104) );
  OAI211X1 U64 ( .A0(n2), .A1(n89), .B0(n88), .C0(n87), .Y(dout[2]) );
  AOI33XL U65 ( .A0(n5), .A1(n98), .A2(n10), .B0(n3), .B1(n94), .B2(n12), .Y(
        n88) );
  AOI222XL U66 ( .A0(n7), .A1(n69), .B0(n2), .B1(n86), .C0(n91), .C1(n14), .Y(
        n87) );
  OAI211X1 U67 ( .A0(n78), .A1(n69), .B0(n77), .C0(n76), .Y(dout[1]) );
  AOI221XL U68 ( .A0(n5), .A1(addr[1]), .B0(n14), .B1(n8), .C0(n72), .Y(n78)
         );
  OAI211X1 U69 ( .A0(n121), .A1(n120), .B0(n119), .C0(n118), .Y(dout[4]) );
  AOI32XL U70 ( .A0(n8), .A1(n114), .A2(addr[5]), .B0(n2), .B1(n112), .Y(n119)
         );
  AOI2BB2X1 U71 ( .B0(n7), .B1(n69), .A0N(n2), .A1N(n117), .Y(n118) );
  BUFX4 U72 ( .A(addr[2]), .Y(n3) );
  CLKINVX3 U73 ( .A(n3), .Y(n6) );
  CLKINVX3 U74 ( .A(n97), .Y(n8) );
endmodule


module sbox6_15 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147;

  NAND2X2 U39 ( .A(n138), .B(addr[3]), .Y(n147) );
  NOR2X2 U47 ( .A(n84), .B(n82), .Y(n138) );
  NOR2X2 U50 ( .A(n14), .B(n4), .Y(n119) );
  NOR2X2 U58 ( .A(n9), .B(n14), .Y(n125) );
  NAND2X2 U61 ( .A(n97), .B(n103), .Y(n112) );
  NOR2X2 U62 ( .A(n18), .B(addr[1]), .Y(n103) );
  NOR2X2 U63 ( .A(n9), .B(addr[3]), .Y(n97) );
  NAND2X2 U64 ( .A(n117), .B(n131), .Y(n140) );
  NOR2X2 U65 ( .A(n5), .B(addr[3]), .Y(n131) );
  NOR2X2 U66 ( .A(n85), .B(addr[6]), .Y(n117) );
  NOR2X1 U1 ( .A(n84), .B(addr[3]), .Y(n102) );
  OAI222X1 U2 ( .A0(n91), .A1(n13), .B0(n3), .B1(n8), .C0(addr[5]), .C1(n10), 
        .Y(n92) );
  CLKINVX1 U3 ( .A(addr[3]), .Y(n1) );
  INVX3 U4 ( .A(addr[3]), .Y(n14) );
  CLKINVX1 U5 ( .A(n9), .Y(n2) );
  INVX4 U6 ( .A(n4), .Y(n9) );
  CLKBUFX3 U7 ( .A(addr[4]), .Y(n4) );
  OAI221X1 U8 ( .A0(n18), .A1(n7), .B0(n14), .B1(n16), .C0(n86), .Y(n90) );
  INVX2 U9 ( .A(n96), .Y(n16) );
  CLKINVX1 U10 ( .A(n84), .Y(n3) );
  BUFX4 U11 ( .A(addr[2]), .Y(n5) );
  NOR2X4 U12 ( .A(addr[1]), .B(addr[6]), .Y(n130) );
  OAI22X1 U13 ( .A0(n14), .A1(n18), .B0(addr[1]), .B1(n10), .Y(n142) );
  OAI221X4 U14 ( .A0(n123), .A1(n17), .B0(n82), .B1(n13), .C0(n15), .Y(n124)
         );
  NOR2X4 U15 ( .A(n5), .B(addr[5]), .Y(n143) );
  INVX1 U16 ( .A(n130), .Y(n83) );
  CLKINVX1 U17 ( .A(n125), .Y(n7) );
  NAND2X1 U18 ( .A(n83), .B(n16), .Y(n105) );
  INVXL U19 ( .A(n121), .Y(n12) );
  CLKINVX1 U20 ( .A(n138), .Y(n81) );
  AOI211X1 U21 ( .A0(n13), .A1(n14), .B0(n131), .C0(n143), .Y(n121) );
  CLKINVX1 U22 ( .A(n117), .Y(n82) );
  CLKINVX1 U23 ( .A(n119), .Y(n10) );
  NOR2X1 U24 ( .A(n16), .B(n123), .Y(n144) );
  NOR2X1 U25 ( .A(n85), .B(n18), .Y(n96) );
  CLKINVX1 U26 ( .A(n103), .Y(n17) );
  OAI211X1 U27 ( .A0(n83), .A1(n7), .B0(n104), .C0(n112), .Y(n108) );
  OAI21XL U28 ( .A0(n103), .A1(n117), .B0(n102), .Y(n104) );
  OAI21XL U29 ( .A0(n132), .A1(n18), .B0(n1), .Y(n86) );
  AOI21X1 U30 ( .A0(n9), .A1(n102), .B0(n125), .Y(n91) );
  OAI2BB2XL U31 ( .B0(n143), .B1(n83), .A0N(n143), .A1N(n117), .Y(n118) );
  CLKINVX1 U32 ( .A(n122), .Y(n15) );
  CLKINVX1 U33 ( .A(n126), .Y(n11) );
  CLKINVX1 U34 ( .A(n97), .Y(n8) );
  NAND2BX1 U35 ( .AN(n144), .B(n137), .Y(n107) );
  CLKINVX1 U36 ( .A(addr[1]), .Y(n85) );
  NOR2X1 U37 ( .A(n16), .B(n3), .Y(n122) );
  NOR2X1 U38 ( .A(addr[1]), .B(n2), .Y(n132) );
  OAI22X1 U40 ( .A0(n10), .A1(n82), .B0(n5), .B1(n11), .Y(n88) );
  NAND2X1 U41 ( .A(n5), .B(n13), .Y(n123) );
  NAND4X1 U42 ( .A(n147), .B(n140), .C(n100), .D(n99), .Y(n101) );
  AOI222XL U43 ( .A0(n98), .A1(n84), .B0(n102), .B1(n130), .C0(n97), .C1(n105), 
        .Y(n99) );
  NAND3X1 U44 ( .A(n5), .B(n10), .C(n96), .Y(n100) );
  OAI221X1 U45 ( .A0(n14), .A1(n17), .B0(n10), .B1(n18), .C0(n11), .Y(n98) );
  AOI22X1 U46 ( .A0(n4), .A1(n115), .B0(addr[5]), .B1(n114), .Y(n129) );
  OAI21XL U48 ( .A0(n121), .A1(n83), .B0(n147), .Y(n115) );
  OAI21XL U49 ( .A0(n113), .A1(n84), .B0(n112), .Y(n114) );
  AOI221XL U51 ( .A0(n119), .A1(n85), .B0(n130), .B1(addr[3]), .C0(n111), .Y(
        n113) );
  OAI22XL U52 ( .A0(n82), .A1(n9), .B0(addr[3]), .B1(n16), .Y(n111) );
  AOI211X1 U53 ( .A0(n4), .A1(n135), .B0(n134), .C0(n133), .Y(n136) );
  OA21XL U54 ( .A0(n1), .A1(n3), .B0(n132), .Y(n133) );
  OAI2BB2XL U55 ( .B0(n2), .B1(n15), .A0N(n131), .A1N(n130), .Y(n134) );
  OAI22X1 U56 ( .A0(n5), .A1(n82), .B0(n84), .B1(n16), .Y(n135) );
  CLKINVX3 U57 ( .A(addr[5]), .Y(n13) );
  AOI2BB2X1 U59 ( .B0(n5), .B1(n130), .A0N(n3), .A1N(n17), .Y(n137) );
  NOR2X1 U60 ( .A(n17), .B(n2), .Y(n126) );
  AOI2BB2XL U67 ( .B0(n143), .B1(n90), .A0N(n89), .A1N(n13), .Y(n94) );
  AOI211X1 U68 ( .A0(n122), .A1(n4), .B0(n88), .C0(n87), .Y(n89) );
  OAI32X1 U69 ( .A0(n17), .A1(n14), .A2(n84), .B0(n81), .B1(n8), .Y(n87) );
  NAND3X1 U70 ( .A(n147), .B(n140), .C(n139), .Y(n141) );
  AOI32X1 U71 ( .A0(n5), .A1(n85), .A2(n4), .B0(n138), .B1(n9), .Y(n139) );
  AO22XL U72 ( .A0(n143), .A1(n2), .B0(n116), .B1(n9), .Y(n120) );
  OAI21XL U73 ( .A0(n3), .A1(n13), .B0(n123), .Y(n116) );
  CLKINVX1 U74 ( .A(n106), .Y(n6) );
  AOI32XL U75 ( .A0(n105), .A1(n9), .A2(n1), .B0(addr[1]), .B1(n125), .Y(n106)
         );
  OAI211X1 U76 ( .A0(n9), .A1(n140), .B0(n110), .C0(n109), .Y(dout[2]) );
  AOI222XL U77 ( .A0(n108), .A1(n13), .B0(n143), .B1(n6), .C0(n119), .C1(n107), 
        .Y(n109) );
  AOI2BB2XL U78 ( .B0(addr[5]), .B1(n101), .A0N(n84), .A1N(n112), .Y(n110) );
  OAI211X1 U79 ( .A0(n2), .A1(n147), .B0(n146), .C0(n145), .Y(dout[4]) );
  AOI222XL U80 ( .A0(n144), .A1(n14), .B0(n143), .B1(n142), .C0(n141), .C1(n13), .Y(n145) );
  OA22X1 U81 ( .A0(n7), .A1(n137), .B0(n136), .B1(n13), .Y(n146) );
  NAND3X1 U82 ( .A(n129), .B(n128), .C(n127), .Y(dout[3]) );
  AOI32XL U83 ( .A0(n120), .A1(n14), .A2(addr[1]), .B0(n119), .B1(n118), .Y(
        n128) );
  AOI222XL U84 ( .A0(n144), .A1(n9), .B0(n126), .B1(n12), .C0(n125), .C1(n124), 
        .Y(n127) );
  NAND3BX1 U85 ( .AN(n95), .B(n94), .C(n93), .Y(dout[1]) );
  OAI222X1 U86 ( .A0(n140), .A1(n4), .B0(n112), .B1(n84), .C0(n16), .C1(n91), 
        .Y(n95) );
  AOI32XL U87 ( .A0(addr[1]), .A1(n13), .A2(n125), .B0(n130), .B1(n92), .Y(n93) );
  CLKINVX3 U88 ( .A(addr[6]), .Y(n18) );
  CLKINVX3 U89 ( .A(n5), .Y(n84) );
endmodule


module sbox7_15 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148;

  OAI222X4 U19 ( .A0(n11), .A1(n129), .B0(n4), .B1(n8), .C0(addr[1]), .C1(n21), 
        .Y(n122) );
  OAI33X4 U33 ( .A0(addr[1]), .A1(n4), .A2(n5), .B0(n9), .B1(n85), .B2(n84), 
        .Y(n97) );
  NOR2X2 U44 ( .A(n87), .B(n4), .Y(n116) );
  NOR2X2 U48 ( .A(addr[1]), .B(addr[6]), .Y(n136) );
  NOR2X2 U51 ( .A(n16), .B(n87), .Y(n125) );
  NOR2X2 U52 ( .A(n9), .B(addr[3]), .Y(n131) );
  NOR2X2 U58 ( .A(n93), .B(n124), .Y(n142) );
  NOR2X2 U60 ( .A(n10), .B(addr[1]), .Y(n93) );
  NOR2X2 U62 ( .A(n83), .B(n3), .Y(n137) );
  NOR2X2 U65 ( .A(n10), .B(n86), .Y(n140) );
  NAND2X1 U1 ( .A(n3), .B(n4), .Y(n119) );
  CLKBUFX3 U2 ( .A(addr[4]), .Y(n4) );
  CLKINVX1 U3 ( .A(n83), .Y(n1) );
  CLKINVX1 U4 ( .A(n85), .Y(n2) );
  CLKBUFX3 U5 ( .A(addr[2]), .Y(n5) );
  OAI31X1 U6 ( .A0(n87), .A1(n83), .A2(n86), .B0(n117), .Y(n121) );
  NOR2X4 U7 ( .A(n86), .B(addr[6]), .Y(n124) );
  OAI22X1 U8 ( .A0(addr[1]), .A1(n21), .B0(n5), .B1(n113), .Y(n100) );
  OAI22X1 U9 ( .A0(n4), .A1(n16), .B0(addr[3]), .B1(n19), .Y(n103) );
  AOI211XL U10 ( .A0(n5), .A1(n7), .B0(n131), .C0(n130), .Y(n132) );
  NOR3XL U11 ( .A(n11), .B(addr[3]), .C(n2), .Y(n130) );
  OAI21XL U12 ( .A0(n3), .A1(n1), .B0(n119), .Y(n89) );
  BUFX4 U13 ( .A(addr[5]), .Y(n3) );
  AOI221XL U14 ( .A0(n140), .A1(n89), .B0(n109), .B1(n7), .C0(n88), .Y(n96) );
  CLKINVX1 U15 ( .A(n140), .Y(n9) );
  OAI2BB2XL U16 ( .B0(n142), .B1(n19), .A0N(n141), .A1N(n140), .Y(n143) );
  CLKINVX1 U17 ( .A(n125), .Y(n14) );
  CLKINVX1 U18 ( .A(n142), .Y(n7) );
  NAND2X1 U20 ( .A(n14), .B(n20), .Y(n105) );
  CLKINVX1 U21 ( .A(n123), .Y(n15) );
  CLKINVX1 U22 ( .A(n109), .Y(n18) );
  NAND2X1 U23 ( .A(n124), .B(n87), .Y(n113) );
  CLKINVX1 U24 ( .A(n137), .Y(n19) );
  NOR2X1 U25 ( .A(n19), .B(n87), .Y(n109) );
  CLKINVX1 U26 ( .A(n136), .Y(n11) );
  OAI22XL U27 ( .A0(n137), .A1(n8), .B0(n86), .B1(n18), .Y(n146) );
  OAI21X1 U28 ( .A0(n83), .A1(n14), .B0(n129), .Y(n141) );
  NAND2X1 U29 ( .A(n116), .B(n16), .Y(n129) );
  CLKINVX1 U30 ( .A(n93), .Y(n6) );
  OAI21XL U31 ( .A0(n119), .A1(n6), .B0(n118), .Y(n120) );
  OAI21XL U32 ( .A0(n125), .A1(n137), .B0(n124), .Y(n118) );
  NOR2X1 U34 ( .A(n16), .B(n21), .Y(n123) );
  CLKINVX1 U35 ( .A(n145), .Y(n21) );
  OAI22XL U36 ( .A0(n137), .A1(n113), .B0(n10), .B1(n15), .Y(n88) );
  CLKINVX1 U37 ( .A(n116), .Y(n84) );
  CLKINVX1 U38 ( .A(n131), .Y(n8) );
  CLKINVX1 U39 ( .A(n134), .Y(n20) );
  NOR2XL U40 ( .A(n125), .B(n83), .Y(n110) );
  CLKINVX1 U41 ( .A(n119), .Y(n17) );
  CLKINVX1 U42 ( .A(n103), .Y(n12) );
  OA21XL U43 ( .A0(n13), .A1(n6), .B0(n117), .Y(n102) );
  CLKINVX1 U45 ( .A(n105), .Y(n13) );
  OAI2BB1XL U46 ( .A0N(n103), .A1N(n124), .B0(n102), .Y(n104) );
  OAI22X1 U47 ( .A0(n16), .A1(n84), .B0(n4), .B1(n20), .Y(n112) );
  NOR4X1 U49 ( .A(n4), .B(addr[3]), .C(n86), .D(n85), .Y(n99) );
  XNOR2X1 U50 ( .A(addr[6]), .B(n5), .Y(n101) );
  AOI211X1 U53 ( .A0(n116), .A1(addr[6]), .B0(n115), .C0(n114), .Y(n128) );
  OAI222X1 U54 ( .A0(n111), .A1(n9), .B0(n110), .B1(n6), .C0(n11), .C1(n18), 
        .Y(n115) );
  OAI2BB2XL U55 ( .B0(n17), .B1(n113), .A0N(n86), .A1N(n112), .Y(n114) );
  OA21XL U56 ( .A0(n87), .A1(n3), .B0(n15), .Y(n111) );
  NAND2X1 U57 ( .A(n5), .B(n136), .Y(n133) );
  CLKINVX1 U59 ( .A(addr[6]), .Y(n10) );
  AOI211X1 U61 ( .A0(n131), .A1(n3), .B0(n92), .C0(n91), .Y(n95) );
  OAI221X1 U63 ( .A0(n86), .A1(n21), .B0(n9), .B1(n19), .C0(n102), .Y(n92) );
  OAI31X1 U64 ( .A0(n87), .A1(n83), .A2(n11), .B0(n90), .Y(n91) );
  AO21XL U66 ( .A0(n119), .A1(n129), .B0(addr[6]), .Y(n90) );
  NOR2X1 U67 ( .A(n83), .B(addr[3]), .Y(n145) );
  AOI21XL U68 ( .A0(addr[3]), .A1(n98), .B0(n97), .Y(n108) );
  OAI2BB1XL U69 ( .A0N(n85), .A1N(n124), .B0(n133), .Y(n98) );
  NAND3X1 U70 ( .A(n136), .B(n87), .C(n3), .Y(n117) );
  NOR2X1 U71 ( .A(addr[3]), .B(n3), .Y(n134) );
  OAI21X1 U72 ( .A0(n5), .A1(n142), .B0(n133), .Y(n138) );
  OAI22XL U73 ( .A0(n142), .A1(n84), .B0(n1), .B1(n132), .Y(n135) );
  AO21X1 U74 ( .A0(n139), .A1(n16), .B0(n138), .Y(n144) );
  OAI21XL U75 ( .A0(n2), .A1(n86), .B0(n6), .Y(n139) );
  OAI221X1 U76 ( .A0(n96), .A1(n85), .B0(n5), .B1(n95), .C0(n94), .Y(dout[1])
         );
  AOI2BB2X1 U77 ( .B0(n93), .B1(n112), .A0N(n133), .A1N(n12), .Y(n94) );
  OAI211X1 U78 ( .A0(n128), .A1(n85), .B0(n127), .C0(n126), .Y(dout[3]) );
  AOI32XL U79 ( .A0(n125), .A1(n1), .A2(n124), .B0(n123), .B1(n136), .Y(n126)
         );
  OAI31X1 U80 ( .A0(n122), .A1(n121), .A2(n120), .B0(n85), .Y(n127) );
  OAI221X1 U81 ( .A0(n3), .A1(n108), .B0(n107), .B1(n16), .C0(n106), .Y(
        dout[2]) );
  AOI32XL U82 ( .A0(n105), .A1(n85), .A2(n140), .B0(n2), .B1(n104), .Y(n106)
         );
  AOI211X1 U83 ( .A0(n101), .A1(n4), .B0(n100), .C0(n99), .Y(n107) );
  NAND2X1 U84 ( .A(n148), .B(n147), .Y(dout[4]) );
  AOI222XL U85 ( .A0(n136), .A1(n141), .B0(n3), .B1(n135), .C0(n134), .C1(n138), .Y(n148) );
  AOI222XL U86 ( .A0(n5), .A1(n146), .B0(n145), .B1(n144), .C0(n143), .C1(n85), 
        .Y(n147) );
  CLKINVX3 U87 ( .A(n3), .Y(n16) );
  CLKINVX3 U88 ( .A(n4), .Y(n83) );
  CLKINVX3 U89 ( .A(n5), .Y(n85) );
  CLKINVX3 U90 ( .A(addr[1]), .Y(n86) );
  CLKINVX3 U91 ( .A(addr[3]), .Y(n87) );
endmodule


module sbox8_15 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132;

  NAND2X2 U41 ( .A(addr[6]), .B(n75), .Y(n131) );
  NAND2X2 U48 ( .A(addr[4]), .B(n9), .Y(n123) );
  NAND2X2 U49 ( .A(n2), .B(n12), .Y(n87) );
  NAND2X2 U50 ( .A(addr[1]), .B(n15), .Y(n124) );
  NAND2X2 U54 ( .A(addr[2]), .B(n6), .Y(n116) );
  NAND2X2 U60 ( .A(addr[6]), .B(addr[1]), .Y(n105) );
  NAND2X2 U61 ( .A(n75), .B(n15), .Y(n108) );
  OAI32X1 U1 ( .A0(n15), .A1(addr[4]), .A2(n92), .B0(n115), .B1(n108), .Y(n96)
         );
  OAI31X1 U2 ( .A0(n123), .A1(addr[6]), .A2(n116), .B0(n109), .Y(n110) );
  AOI222X1 U3 ( .A0(n88), .A1(addr[2]), .B0(n12), .B1(n7), .C0(n10), .C1(n92), 
        .Y(n114) );
  OAI222X1 U4 ( .A0(addr[2]), .A1(n126), .B0(n9), .B1(n125), .C0(n124), .C1(
        n123), .Y(n127) );
  OAI221X1 U5 ( .A0(n105), .A1(n87), .B0(addr[4]), .B1(n108), .C0(n86), .Y(n90) );
  NAND2X4 U6 ( .A(addr[4]), .B(n2), .Y(n115) );
  AOI32XL U7 ( .A0(n13), .A1(n5), .A2(n2), .B0(n14), .B1(n117), .Y(n130) );
  OA21XL U8 ( .A0(n10), .A1(n6), .B0(n121), .Y(n78) );
  INVXL U9 ( .A(n119), .Y(n3) );
  INVX3 U10 ( .A(n2), .Y(n9) );
  BUFX4 U11 ( .A(addr[3]), .Y(n2) );
  CLKBUFX3 U12 ( .A(addr[5]), .Y(n1) );
  CLKINVX1 U13 ( .A(n108), .Y(n14) );
  CLKINVX1 U14 ( .A(n107), .Y(n4) );
  CLKINVX1 U15 ( .A(n93), .Y(n8) );
  NAND2X1 U16 ( .A(n9), .B(n12), .Y(n93) );
  NAND2X1 U17 ( .A(n10), .B(n6), .Y(n121) );
  OAI21XL U18 ( .A0(n115), .A1(n6), .B0(n107), .Y(n77) );
  OAI21X1 U19 ( .A0(n12), .A1(n6), .B0(n123), .Y(n88) );
  OAI31XL U20 ( .A0(n115), .A1(n75), .A2(n116), .B0(n118), .Y(n94) );
  CLKINVX1 U21 ( .A(n131), .Y(n74) );
  NAND2X1 U22 ( .A(n5), .B(n9), .Y(n107) );
  OAI22XL U23 ( .A0(n116), .A1(n123), .B0(n5), .B1(n115), .Y(n117) );
  OAI22XL U24 ( .A0(n123), .A1(n108), .B0(n131), .B1(n93), .Y(n95) );
  OAI2BB2XL U25 ( .B0(n115), .B1(n131), .A0N(n88), .A1N(n16), .Y(n89) );
  AOI211XL U26 ( .A0(n108), .A1(n105), .B0(n12), .C0(n121), .Y(n85) );
  CLKINVX1 U27 ( .A(n124), .Y(n13) );
  OAI22XL U28 ( .A0(n5), .A1(n123), .B0(n78), .B1(n87), .Y(n81) );
  NAND2BX2 U29 ( .AN(n78), .B(n9), .Y(n120) );
  NAND2XL U30 ( .A(n115), .B(n93), .Y(n104) );
  OAI2BB2XL U31 ( .B0(n106), .B1(n105), .A0N(n104), .A1N(n13), .Y(n111) );
  NOR2BXL U32 ( .AN(n123), .B(n103), .Y(n106) );
  NAND3X1 U33 ( .A(n104), .B(n75), .C(n5), .Y(n84) );
  AO21X1 U34 ( .A0(n5), .A1(n16), .B0(n101), .Y(n102) );
  OAI33X1 U35 ( .A0(n15), .A1(n9), .A2(n100), .B0(n10), .B1(n103), .B2(n124), 
        .Y(n101) );
  OA22XL U36 ( .A0(n107), .A1(n131), .B0(n120), .B1(n124), .Y(n98) );
  CLKINVX1 U37 ( .A(n125), .Y(n11) );
  OAI21XL U38 ( .A0(n13), .A1(n74), .B0(addr[4]), .Y(n86) );
  NAND2X1 U39 ( .A(n1), .B(n10), .Y(n100) );
  OAI221X1 U40 ( .A0(n124), .A1(n121), .B0(addr[1]), .B1(n120), .C0(n3), .Y(
        n128) );
  OAI31XL U42 ( .A0(n10), .A1(n75), .A2(n9), .B0(n118), .Y(n119) );
  NAND2X1 U43 ( .A(n16), .B(addr[2]), .Y(n125) );
  NAND4XL U44 ( .A(n74), .B(n1), .C(n2), .D(addr[2]), .Y(n109) );
  NAND3X1 U45 ( .A(n5), .B(n15), .C(n2), .Y(n118) );
  OAI21XL U46 ( .A0(n1), .A1(n87), .B0(n114), .Y(n76) );
  OAI22XL U47 ( .A0(n108), .A1(n120), .B0(n79), .B1(n100), .Y(n80) );
  AOI221XL U51 ( .A0(n74), .A1(n9), .B0(n16), .B1(n2), .C0(n91), .Y(n79) );
  NOR2X1 U52 ( .A(n1), .B(n2), .Y(n103) );
  NOR2X1 U53 ( .A(n87), .B(addr[6]), .Y(n91) );
  NOR2X1 U55 ( .A(n9), .B(n1), .Y(n92) );
  CLKINVX1 U56 ( .A(n100), .Y(n7) );
  OA21XL U57 ( .A0(n1), .A1(n115), .B0(n120), .Y(n132) );
  AOI221XL U58 ( .A0(n14), .A1(n2), .B0(n16), .B1(addr[4]), .C0(n122), .Y(n126) );
  OAI22XL U59 ( .A0(n2), .A1(n75), .B0(addr[4]), .B1(n131), .Y(n122) );
  OAI211X1 U62 ( .A0(addr[2]), .A1(n99), .B0(n98), .C0(n97), .Y(dout[2]) );
  AOI221XL U63 ( .A0(addr[2]), .A1(n96), .B0(n1), .B1(n95), .C0(n94), .Y(n97)
         );
  AOI221XL U64 ( .A0(n91), .A1(n1), .B0(n90), .B1(n6), .C0(n89), .Y(n99) );
  OAI211X1 U65 ( .A0(n132), .A1(n131), .B0(n130), .C0(n129), .Y(dout[4]) );
  AOI222XL U66 ( .A0(n128), .A1(n12), .B0(n1), .B1(n127), .C0(n4), .C1(n16), 
        .Y(n129) );
  OAI211X1 U67 ( .A0(addr[1]), .A1(n114), .B0(n113), .C0(n112), .Y(dout[3]) );
  AOI221XL U68 ( .A0(n111), .A1(n10), .B0(n4), .B1(n14), .C0(n110), .Y(n112)
         );
  AOI2BB2XL U69 ( .B0(n102), .B1(n12), .A0N(n115), .A1N(n125), .Y(n113) );
  NAND4BX1 U70 ( .AN(n85), .B(n84), .C(n83), .D(n82), .Y(dout[1]) );
  AOI221XL U71 ( .A0(n74), .A1(n81), .B0(n8), .B1(n11), .C0(n80), .Y(n82) );
  AOI22X1 U72 ( .A0(n16), .A1(n77), .B0(n13), .B1(n76), .Y(n83) );
  CLKINVX3 U73 ( .A(n116), .Y(n5) );
  CLKINVX3 U74 ( .A(n1), .Y(n6) );
  CLKINVX3 U75 ( .A(addr[2]), .Y(n10) );
  CLKINVX3 U76 ( .A(addr[4]), .Y(n12) );
  CLKINVX3 U77 ( .A(addr[6]), .Y(n15) );
  CLKINVX3 U78 ( .A(n105), .Y(n16) );
  CLKINVX3 U79 ( .A(addr[1]), .Y(n75) );
endmodule


module crp_15 ( P, R, K_sub );
  output [1:32] P;
  input [1:32] R;
  input [1:48] K_sub;
  wire   n1;
  wire   [1:48] X;

  sbox1_15 u0 ( .addr(X[1:6]), .dout({P[9], P[17], P[23], P[31]}) );
  sbox2_15 u1 ( .addr({X[7], n1, X[9:12]}), .dout({P[13], P[28], P[2], P[18]})
         );
  sbox3_15 u2 ( .addr(X[13:18]), .dout({P[24], P[16], P[30], P[6]}) );
  sbox4_15 u3 ( .addr(X[19:24]), .dout({P[26], P[20], P[10], P[1]}) );
  sbox5_15 u4 ( .addr(X[25:30]), .dout({P[8], P[14], P[25], P[3]}) );
  sbox6_15 u5 ( .addr(X[31:36]), .dout({P[4], P[29], P[11], P[19]}) );
  sbox7_15 u6 ( .addr(X[37:42]), .dout({P[32], P[12], P[22], P[7]}) );
  sbox8_15 u7 ( .addr(X[43:48]), .dout({P[5], P[27], P[15], P[21]}) );
  XNOR2X1 U1 ( .A(R[5]), .B(K_sub[8]), .Y(X[8]) );
  INVX3 U2 ( .A(X[8]), .Y(n1) );
  XOR2X1 U3 ( .A(R[1]), .B(K_sub[2]), .Y(X[2]) );
  CLKXOR2X4 U4 ( .A(R[29]), .B(K_sub[42]), .Y(X[42]) );
  CLKXOR2X4 U5 ( .A(R[16]), .B(K_sub[25]), .Y(X[25]) );
  CLKXOR2X4 U6 ( .A(R[8]), .B(K_sub[11]), .Y(X[11]) );
  CLKXOR2X4 U7 ( .A(R[20]), .B(K_sub[31]), .Y(X[31]) );
  CLKXOR2X4 U8 ( .A(R[29]), .B(K_sub[44]), .Y(X[44]) );
  CLKXOR2X4 U9 ( .A(R[16]), .B(K_sub[23]), .Y(X[23]) );
  CLKXOR2X4 U10 ( .A(R[10]), .B(K_sub[15]), .Y(X[15]) );
  CLKXOR2X4 U11 ( .A(R[31]), .B(K_sub[46]), .Y(X[46]) );
  CLKXOR2X4 U12 ( .A(R[22]), .B(K_sub[33]), .Y(X[33]) );
  CLKXOR2X4 U13 ( .A(R[12]), .B(K_sub[19]), .Y(X[19]) );
  CLKXOR2X4 U14 ( .A(R[26]), .B(K_sub[39]), .Y(X[39]) );
  CLKXOR2X4 U15 ( .A(R[20]), .B(K_sub[29]), .Y(X[29]) );
  CLKXOR2X2 U16 ( .A(R[4]), .B(K_sub[5]), .Y(X[5]) );
  CLKXOR2X2 U17 ( .A(R[15]), .B(K_sub[22]), .Y(X[22]) );
  CLKXOR2X2 U18 ( .A(R[24]), .B(K_sub[35]), .Y(X[35]) );
  CLKXOR2X2 U19 ( .A(R[21]), .B(K_sub[30]), .Y(X[30]) );
  CLKXOR2X2 U20 ( .A(R[12]), .B(K_sub[17]), .Y(X[17]) );
  CLKXOR2X2 U21 ( .A(R[32]), .B(K_sub[1]), .Y(X[1]) );
  CLKXOR2X2 U22 ( .A(R[13]), .B(K_sub[20]), .Y(X[20]) );
  CLKXOR2X2 U23 ( .A(R[18]), .B(K_sub[27]), .Y(X[27]) );
  CLKXOR2X2 U24 ( .A(R[8]), .B(K_sub[13]), .Y(X[13]) );
  CLKXOR2X2 U25 ( .A(R[5]), .B(K_sub[6]), .Y(X[6]) );
  CLKXOR2X2 U26 ( .A(R[4]), .B(K_sub[7]), .Y(X[7]) );
  CLKXOR2X2 U27 ( .A(R[24]), .B(K_sub[37]), .Y(X[37]) );
  CLKXOR2X2 U28 ( .A(R[28]), .B(K_sub[43]), .Y(X[43]) );
  CLKXOR2X2 U29 ( .A(R[1]), .B(K_sub[48]), .Y(X[48]) );
  CLKXOR2X2 U30 ( .A(R[17]), .B(K_sub[24]), .Y(X[24]) );
  CLKXOR2X2 U31 ( .A(R[9]), .B(K_sub[12]), .Y(X[12]) );
  CLKXOR2X2 U32 ( .A(R[13]), .B(K_sub[18]), .Y(X[18]) );
  CLKXOR2X2 U33 ( .A(R[25]), .B(K_sub[36]), .Y(X[36]) );
  XOR2X1 U34 ( .A(R[23]), .B(K_sub[34]), .Y(X[34]) );
  XOR2X1 U35 ( .A(R[9]), .B(K_sub[14]), .Y(X[14]) );
  XOR2X1 U36 ( .A(R[30]), .B(K_sub[45]), .Y(X[45]) );
  XOR2X1 U37 ( .A(R[21]), .B(K_sub[32]), .Y(X[32]) );
  XOR2X1 U38 ( .A(R[25]), .B(K_sub[38]), .Y(X[38]) );
  XOR2X1 U39 ( .A(R[27]), .B(K_sub[40]), .Y(X[40]) );
  XOR2X1 U40 ( .A(R[3]), .B(K_sub[4]), .Y(X[4]) );
  XOR2X1 U41 ( .A(R[11]), .B(K_sub[16]), .Y(X[16]) );
  XOR2X1 U42 ( .A(R[7]), .B(K_sub[10]), .Y(X[10]) );
  XOR2X1 U43 ( .A(R[14]), .B(K_sub[21]), .Y(X[21]) );
  XOR2X1 U44 ( .A(R[6]), .B(K_sub[9]), .Y(X[9]) );
  XOR2X1 U45 ( .A(R[2]), .B(K_sub[3]), .Y(X[3]) );
  XOR2X1 U46 ( .A(R[28]), .B(K_sub[41]), .Y(X[41]) );
  XOR2X1 U47 ( .A(R[17]), .B(K_sub[26]), .Y(X[26]) );
  XOR2X1 U48 ( .A(R[32]), .B(K_sub[47]), .Y(X[47]) );
  XOR2X1 U49 ( .A(R[19]), .B(K_sub[28]), .Y(X[28]) );
endmodule


module sbox1_14 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127;

  OAI222X4 U13 ( .A0(addr[5]), .A1(n101), .B0(n1), .B1(n100), .C0(n99), .C1(n9), .Y(dout[3]) );
  OAI21X2 U42 ( .A0(n4), .A1(n112), .B0(n106), .Y(n123) );
  NAND2X2 U44 ( .A(addr[6]), .B(n69), .Y(n115) );
  NAND2X2 U48 ( .A(addr[1]), .B(n72), .Y(n114) );
  OAI22X2 U49 ( .A0(n11), .A1(n10), .B0(addr[5]), .B1(n120), .Y(n85) );
  NAND2X2 U50 ( .A(n3), .B(n11), .Y(n120) );
  NOR2X2 U51 ( .A(n11), .B(n3), .Y(n124) );
  NOR3X2 U55 ( .A(n2), .B(addr[6]), .C(n9), .Y(n102) );
  NOR2X2 U56 ( .A(n109), .B(n3), .Y(n93) );
  NAND2X2 U57 ( .A(addr[1]), .B(addr[6]), .Y(n109) );
  NAND2X2 U59 ( .A(n69), .B(n72), .Y(n112) );
  NOR2X1 U1 ( .A(n114), .B(n120), .Y(n104) );
  BUFX4 U2 ( .A(addr[4]), .Y(n2) );
  CLKBUFX3 U3 ( .A(addr[2]), .Y(n1) );
  OAI32X1 U4 ( .A0(n112), .A1(n2), .A2(n4), .B0(n115), .B1(n113), .Y(n80) );
  NOR2BXL U5 ( .AN(n118), .B(n1), .Y(n122) );
  CLKBUFX3 U6 ( .A(addr[2]), .Y(n4) );
  INVX3 U7 ( .A(addr[6]), .Y(n72) );
  OAI221X4 U8 ( .A0(n88), .A1(n10), .B0(addr[5]), .B1(n87), .C0(n86), .Y(
        dout[2]) );
  OAI221X4 U9 ( .A0(addr[5]), .A1(n127), .B0(n126), .B1(n10), .C0(n125), .Y(
        dout[4]) );
  OA21XL U10 ( .A0(n95), .A1(n115), .B0(n107), .Y(n119) );
  AOI222XL U11 ( .A0(n13), .A1(n1), .B0(n2), .B1(n110), .C0(n70), .C1(n9), .Y(
        n111) );
  AOI2BB2X1 U12 ( .B0(n2), .B1(n70), .A0N(addr[4]), .A1N(n115), .Y(n91) );
  BUFX4 U14 ( .A(addr[3]), .Y(n3) );
  CLKINVX1 U15 ( .A(n112), .Y(n13) );
  CLKINVX1 U16 ( .A(n113), .Y(n5) );
  NAND2BX1 U17 ( .AN(n104), .B(n119), .Y(n84) );
  CLKXOR2X2 U18 ( .A(n6), .B(n9), .Y(n90) );
  NOR2X1 U19 ( .A(n11), .B(n6), .Y(n118) );
  OAI21XL U20 ( .A0(n6), .A1(n114), .B0(n91), .Y(n92) );
  NAND2X1 U21 ( .A(n93), .B(n11), .Y(n107) );
  NAND2X1 U22 ( .A(n9), .B(n6), .Y(n113) );
  OAI211X1 U23 ( .A0(n11), .A1(n114), .B0(n108), .C0(n107), .Y(n89) );
  CLKINVX1 U24 ( .A(n109), .Y(n70) );
  NAND2X1 U25 ( .A(n124), .B(n12), .Y(n108) );
  CLKINVX1 U26 ( .A(n114), .Y(n71) );
  CLKINVX1 U27 ( .A(n115), .Y(n12) );
  CLKINVX1 U28 ( .A(n95), .Y(n8) );
  AO22X1 U29 ( .A0(n90), .A1(n12), .B0(n6), .B1(n123), .Y(n76) );
  OAI31X1 U30 ( .A0(n9), .A1(n3), .A2(n69), .B0(n103), .Y(n105) );
  AOI31XL U31 ( .A0(n69), .A1(n9), .A2(n2), .B0(n102), .Y(n103) );
  AOI211X1 U32 ( .A0(n7), .A1(n4), .B0(n117), .C0(n116), .Y(n126) );
  CLKINVX1 U33 ( .A(n108), .Y(n7) );
  AOI211X1 U34 ( .A0(n115), .A1(n114), .B0(n113), .C0(n2), .Y(n116) );
  OAI22X1 U35 ( .A0(n120), .A1(n112), .B0(n111), .B1(n6), .Y(n117) );
  AOI211X1 U36 ( .A0(n70), .A1(n118), .B0(n81), .C0(n80), .Y(n88) );
  OAI22X1 U37 ( .A0(n91), .A1(n9), .B0(n3), .B1(n106), .Y(n81) );
  CLKINVX3 U38 ( .A(addr[5]), .Y(n10) );
  NAND2X1 U39 ( .A(n3), .B(n10), .Y(n95) );
  NAND2X1 U40 ( .A(n71), .B(n1), .Y(n106) );
  XOR2X1 U41 ( .A(n82), .B(n2), .Y(n83) );
  NAND2X1 U43 ( .A(n1), .B(n3), .Y(n82) );
  OAI22XL U45 ( .A0(n3), .A1(n69), .B0(n6), .B1(n112), .Y(n94) );
  AOI211XL U46 ( .A0(n98), .A1(n6), .B0(n97), .C0(n104), .Y(n99) );
  OAI22XL U47 ( .A0(n96), .A1(n11), .B0(n95), .B1(n109), .Y(n97) );
  OAI22XL U52 ( .A0(n72), .A1(n10), .B0(n2), .B1(addr[1]), .Y(n98) );
  AOI221XL U53 ( .A0(n8), .A1(addr[6]), .B0(addr[5]), .B1(n94), .C0(n93), .Y(
        n96) );
  OAI21XL U54 ( .A0(addr[1]), .A1(n120), .B0(n119), .Y(n121) );
  AOI221XL U58 ( .A0(n13), .A1(n118), .B0(n93), .B1(n10), .C0(n75), .Y(n78) );
  OAI31X1 U60 ( .A0(n10), .A1(n2), .A2(n74), .B0(n73), .Y(n75) );
  OA21XL U61 ( .A0(n3), .A1(n72), .B0(n109), .Y(n74) );
  OAI21XL U62 ( .A0(n124), .A1(n85), .B0(n71), .Y(n73) );
  OAI21XL U63 ( .A0(n1), .A1(n69), .B0(n109), .Y(n110) );
  INVX4 U64 ( .A(n4), .Y(n9) );
  AOI222XL U65 ( .A0(n124), .A1(n123), .B0(n122), .B1(addr[6]), .C0(n1), .C1(
        n121), .Y(n125) );
  NOR4BBX1 U66 ( .AN(n107), .BN(n106), .C(n105), .D(n104), .Y(n127) );
  AOI222XL U67 ( .A0(n13), .A1(n90), .B0(n89), .B1(n9), .C0(n123), .C1(n11), 
        .Y(n101) );
  AOI2BB2XL U68 ( .B0(addr[5]), .B1(n92), .A0N(n120), .A1N(addr[1]), .Y(n100)
         );
  AOI32X1 U69 ( .A0(n4), .A1(n85), .A2(n13), .B0(n84), .B1(n9), .Y(n86) );
  AOI222XL U70 ( .A0(n124), .A1(n69), .B0(n83), .B1(addr[1]), .C0(n5), .C1(n72), .Y(n87) );
  OAI221X1 U71 ( .A0(n79), .A1(n10), .B0(n4), .B1(n78), .C0(n77), .Y(dout[1])
         );
  AOI32XL U72 ( .A0(addr[6]), .A1(n85), .A2(n1), .B0(n76), .B1(n10), .Y(n77)
         );
  AOI221X1 U73 ( .A0(n13), .A1(n90), .B0(n4), .B1(n93), .C0(n102), .Y(n79) );
  CLKINVX3 U74 ( .A(n3), .Y(n6) );
  CLKINVX3 U75 ( .A(n2), .Y(n11) );
  CLKINVX3 U76 ( .A(addr[1]), .Y(n69) );
endmodule


module sbox2_14 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147;

  NAND2X2 U55 ( .A(n2), .B(n16), .Y(n136) );
  NAND2X2 U57 ( .A(addr[2]), .B(n83), .Y(n104) );
  NAND2X2 U60 ( .A(addr[5]), .B(addr[2]), .Y(n132) );
  NOR2X2 U61 ( .A(n7), .B(n4), .Y(n101) );
  NAND2X2 U62 ( .A(n6), .B(n9), .Y(n146) );
  NAND2X2 U63 ( .A(n3), .B(n11), .Y(n124) );
  NAND2X2 U64 ( .A(addr[6]), .B(n6), .Y(n122) );
  NAND2X2 U67 ( .A(n3), .B(n2), .Y(n133) );
  AOI222XL U1 ( .A0(n15), .A1(n8), .B0(n88), .B1(n11), .C0(n140), .C1(n4), .Y(
        n89) );
  CLKINVX1 U2 ( .A(n121), .Y(n7) );
  CLKINVX1 U3 ( .A(addr[5]), .Y(n1) );
  INVX3 U4 ( .A(addr[5]), .Y(n83) );
  OAI211X4 U5 ( .A0(n147), .A1(n146), .B0(n145), .C0(n144), .Y(dout[4]) );
  NOR2X1 U6 ( .A(n104), .B(n2), .Y(n141) );
  NOR2X1 U7 ( .A(n124), .B(n2), .Y(n140) );
  CLKBUFX4 U8 ( .A(addr[4]), .Y(n2) );
  NAND3XL U9 ( .A(n98), .B(n97), .C(n96), .Y(dout[1]) );
  NAND2X1 U10 ( .A(addr[1]), .B(addr[6]), .Y(n121) );
  CLKINVX2 U11 ( .A(addr[1]), .Y(n6) );
  OAI221X1 U12 ( .A0(addr[1]), .A1(n136), .B0(n133), .B1(n6), .C0(n87), .Y(n95) );
  NAND2X4 U13 ( .A(addr[1]), .B(n9), .Y(n114) );
  INVX3 U14 ( .A(addr[6]), .Y(n9) );
  NAND2XL U15 ( .A(n102), .B(n16), .Y(n109) );
  AOI211XL U16 ( .A0(n12), .A1(n95), .B0(n94), .C0(n93), .Y(n96) );
  AOI2BB2X1 U17 ( .B0(n83), .B1(n10), .A0N(n104), .A1N(n136), .Y(n117) );
  NOR3BXL U18 ( .AN(n135), .B(n134), .C(n15), .Y(n147) );
  BUFX4 U19 ( .A(addr[3]), .Y(n3) );
  NAND2X1 U20 ( .A(n15), .B(n7), .Y(n113) );
  CLKINVX1 U21 ( .A(n146), .Y(n4) );
  CLKINVX1 U22 ( .A(n115), .Y(n15) );
  CLKINVX1 U23 ( .A(n122), .Y(n5) );
  OAI31X1 U24 ( .A0(n124), .A1(n9), .A2(n83), .B0(n123), .Y(n128) );
  OAI21XL U25 ( .A0(n83), .A1(n6), .B0(n140), .Y(n123) );
  OAI22X1 U26 ( .A0(n122), .A1(n124), .B0(n101), .B1(n132), .Y(n84) );
  INVX1 U27 ( .A(n114), .Y(n8) );
  OAI22X1 U28 ( .A0(n122), .A1(n16), .B0(n82), .B1(n121), .Y(n129) );
  NAND3X1 U29 ( .A(n82), .B(n83), .C(n6), .Y(n111) );
  NAND2X1 U30 ( .A(n16), .B(n82), .Y(n115) );
  OAI21XL U31 ( .A0(n11), .A1(n133), .B0(n135), .Y(n85) );
  OAI22XL U32 ( .A0(n117), .A1(n146), .B0(n116), .B1(n132), .Y(n118) );
  AOI222XL U33 ( .A0(n8), .A1(n115), .B0(n81), .B1(n9), .C0(n15), .C1(n4), .Y(
        n116) );
  CLKINVX1 U34 ( .A(n104), .Y(n13) );
  OAI2BB2XL U35 ( .B0(n114), .B1(n135), .A0N(n126), .A1N(n81), .Y(n106) );
  OAI21XL U36 ( .A0(n112), .A1(n114), .B0(n111), .Y(n120) );
  OAI21XL U37 ( .A0(n133), .A1(n114), .B0(n113), .Y(n119) );
  CLKINVX1 U38 ( .A(n124), .Y(n10) );
  CLKINVX1 U39 ( .A(n136), .Y(n14) );
  CLKINVX1 U40 ( .A(n133), .Y(n81) );
  CLKINVX1 U41 ( .A(n132), .Y(n12) );
  AOI2BB1X1 U42 ( .A0N(n126), .A1N(n125), .B0(n136), .Y(n127) );
  OAI22XL U43 ( .A0(n104), .A1(n114), .B0(n101), .B1(n132), .Y(n102) );
  AO21XL U44 ( .A0(n11), .A1(n14), .B0(n141), .Y(n86) );
  AO21X1 U45 ( .A0(n16), .A1(n13), .B0(n140), .Y(n142) );
  NAND3X1 U46 ( .A(n11), .B(n82), .C(addr[5]), .Y(n135) );
  OAI22X1 U47 ( .A0(addr[5]), .A1(n121), .B0(n122), .B1(n83), .Y(n126) );
  AOI2BB1X1 U48 ( .A0N(n3), .A1N(n1), .B0(n14), .Y(n112) );
  NOR3X1 U49 ( .A(addr[1]), .B(addr[2]), .C(n83), .Y(n125) );
  AOI2BB1XL U50 ( .A0N(n92), .A1N(n91), .B0(addr[5]), .Y(n93) );
  OAI22XL U51 ( .A0(n117), .A1(n114), .B0(n89), .B1(n1), .Y(n94) );
  OAI31XL U52 ( .A0(n114), .A1(n2), .A2(n16), .B0(n90), .Y(n91) );
  OAI21XL U53 ( .A0(n81), .A1(n10), .B0(n5), .Y(n90) );
  NAND2X1 U54 ( .A(n8), .B(n2), .Y(n137) );
  OAI31XL U56 ( .A0(n101), .A1(n3), .A2(addr[2]), .B0(n113), .Y(n92) );
  OAI211X1 U58 ( .A0(n139), .A1(n83), .B0(n138), .C0(n137), .Y(n143) );
  NAND3X1 U59 ( .A(n82), .B(n83), .C(addr[6]), .Y(n138) );
  AOI2BB2X1 U65 ( .B0(n5), .B1(n16), .A0N(n6), .A1N(n136), .Y(n139) );
  OAI22XL U66 ( .A0(addr[5]), .A1(n133), .B0(n3), .B1(n132), .Y(n134) );
  OAI2BB2XL U68 ( .B0(n112), .B1(n122), .A0N(n1), .A1N(n99), .Y(n100) );
  OAI211X1 U69 ( .A0(n146), .A1(n2), .B0(n137), .C0(n113), .Y(n99) );
  NAND3X1 U70 ( .A(n5), .B(n82), .C(n3), .Y(n87) );
  AOI2BB2XL U71 ( .B0(n3), .B1(n105), .A0N(n137), .A1N(n132), .Y(n108) );
  OAI211XL U72 ( .A0(n104), .A1(n146), .B0(n103), .C0(n111), .Y(n105) );
  NAND3XL U73 ( .A(addr[5]), .B(n82), .C(n7), .Y(n103) );
  OAI22XL U74 ( .A0(n3), .A1(n114), .B0(n9), .B1(n115), .Y(n88) );
  NAND4X1 U75 ( .A(n110), .B(n109), .C(n108), .D(n107), .Y(dout[2]) );
  AOI32XL U76 ( .A0(addr[1]), .A1(addr[2]), .A2(n14), .B0(n100), .B1(n11), .Y(
        n110) );
  AOI221XL U77 ( .A0(n125), .A1(addr[4]), .B0(n141), .B1(n5), .C0(n106), .Y(
        n107) );
  AOI33XL U78 ( .A0(n5), .A1(n13), .A2(n2), .B0(n12), .B1(n146), .B2(n3), .Y(
        n145) );
  AOI222XL U79 ( .A0(n143), .A1(n11), .B0(n7), .B1(n142), .C0(n8), .C1(n141), 
        .Y(n144) );
  AOI32XL U80 ( .A0(n13), .A1(n6), .A2(n15), .B0(n4), .B1(n86), .Y(n97) );
  AOI22X1 U81 ( .A0(n7), .A1(n85), .B0(n2), .B1(n84), .Y(n98) );
  NAND2X1 U82 ( .A(n131), .B(n130), .Y(dout[3]) );
  AOI221XL U83 ( .A0(n120), .A1(n11), .B0(addr[2]), .B1(n119), .C0(n118), .Y(
        n131) );
  AOI211X1 U84 ( .A0(n13), .A1(n129), .B0(n128), .C0(n127), .Y(n130) );
  CLKINVX3 U85 ( .A(addr[2]), .Y(n11) );
  CLKINVX3 U86 ( .A(n3), .Y(n16) );
  CLKINVX3 U87 ( .A(n2), .Y(n82) );
endmodule


module sbox3_14 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134;

  NOR2X2 U35 ( .A(n7), .B(addr[3]), .Y(n109) );
  NOR2X2 U50 ( .A(addr[1]), .B(addr[6]), .Y(n108) );
  NOR2X2 U52 ( .A(n14), .B(n3), .Y(n88) );
  NOR2X2 U56 ( .A(n14), .B(n15), .Y(n95) );
  NOR2X1 U1 ( .A(n7), .B(n14), .Y(n107) );
  OAI221X1 U2 ( .A0(n125), .A1(n7), .B0(n4), .B1(addr[1]), .C0(n78), .Y(n105)
         );
  INVXL U3 ( .A(n2), .Y(n1) );
  NOR2X1 U4 ( .A(n20), .B(n4), .Y(n92) );
  NOR2X1 U5 ( .A(n9), .B(n4), .Y(n122) );
  NOR2X1 U6 ( .A(n78), .B(n4), .Y(n96) );
  CLKBUFX3 U7 ( .A(addr[2]), .Y(n4) );
  INVX1 U8 ( .A(addr[2]), .Y(n2) );
  NOR2X1 U9 ( .A(n4), .B(n3), .Y(n111) );
  BUFX4 U10 ( .A(addr[4]), .Y(n3) );
  OAI33X1 U11 ( .A0(n9), .A1(n126), .A2(n15), .B0(n7), .B1(n95), .B2(n120), 
        .Y(n80) );
  INVX3 U12 ( .A(n4), .Y(n15) );
  OAI221X1 U13 ( .A0(addr[5]), .A1(n91), .B0(n90), .B1(n17), .C0(n89), .Y(
        dout[1]) );
  NOR2X4 U14 ( .A(n76), .B(n79), .Y(n125) );
  NOR2X4 U15 ( .A(addr[3]), .B(n3), .Y(n131) );
  NOR2X4 U16 ( .A(n79), .B(addr[6]), .Y(n126) );
  INVX3 U17 ( .A(addr[1]), .Y(n79) );
  NAND2XL U18 ( .A(n95), .B(n125), .Y(n133) );
  OAI211XL U19 ( .A0(n3), .A1(n16), .B0(n129), .C0(n128), .Y(n130) );
  NAND4XL U20 ( .A(n115), .B(n114), .C(n113), .D(n112), .Y(n116) );
  CLKINVX1 U21 ( .A(n133), .Y(n13) );
  INVX1 U22 ( .A(n125), .Y(n18) );
  CLKINVX1 U23 ( .A(n107), .Y(n5) );
  NAND2X1 U24 ( .A(n20), .B(n6), .Y(n123) );
  CLKINVX1 U25 ( .A(n87), .Y(n6) );
  CLKINVX1 U26 ( .A(n121), .Y(n12) );
  CLKINVX1 U27 ( .A(n120), .Y(n19) );
  CLKINVX1 U28 ( .A(n115), .Y(n10) );
  CLKINVX1 U29 ( .A(n108), .Y(n78) );
  NOR2X1 U30 ( .A(n20), .B(n15), .Y(n104) );
  NOR2X1 U31 ( .A(n18), .B(n15), .Y(n110) );
  INVX1 U32 ( .A(n126), .Y(n77) );
  AOI21X1 U33 ( .A0(n14), .A1(n15), .B0(n95), .Y(n121) );
  OAI21XL U34 ( .A0(n111), .A1(n131), .B0(n125), .Y(n83) );
  CLKINVX1 U36 ( .A(n82), .Y(n20) );
  NOR2X1 U37 ( .A(n77), .B(n7), .Y(n87) );
  NOR2X1 U38 ( .A(n125), .B(n108), .Y(n120) );
  OAI21XL U39 ( .A0(n110), .A1(n92), .B0(n131), .Y(n101) );
  NAND2X1 U40 ( .A(n104), .B(n88), .Y(n115) );
  CLKINVX1 U41 ( .A(n88), .Y(n9) );
  CLKINVX1 U42 ( .A(n92), .Y(n16) );
  CLKINVX1 U43 ( .A(n111), .Y(n11) );
  CLKINVX1 U44 ( .A(n122), .Y(n8) );
  OR2X1 U45 ( .A(n104), .B(n96), .Y(n127) );
  OAI221X1 U46 ( .A0(n77), .A1(n11), .B0(n15), .B1(n6), .C0(n94), .Y(n99) );
  AOI221XL U47 ( .A0(n96), .A1(n3), .B0(n93), .B1(n7), .C0(n13), .Y(n94) );
  OAI21XL U48 ( .A0(n15), .A1(n78), .B0(n16), .Y(n93) );
  XNOR2X1 U49 ( .A(addr[5]), .B(addr[3]), .Y(n103) );
  CLKINVX1 U51 ( .A(addr[5]), .Y(n17) );
  OAI221X1 U53 ( .A0(n78), .A1(n11), .B0(n18), .B1(n9), .C0(n106), .Y(n117) );
  AOI221XL U54 ( .A0(addr[3]), .A1(n105), .B0(n104), .B1(n131), .C0(n13), .Y(
        n106) );
  CLKINVX1 U55 ( .A(addr[6]), .Y(n76) );
  NAND3X1 U57 ( .A(n4), .B(n79), .C(n109), .Y(n114) );
  NOR2X1 U58 ( .A(n76), .B(addr[1]), .Y(n82) );
  AOI32XL U59 ( .A0(n15), .A1(n14), .A2(n125), .B0(n124), .B1(n76), .Y(n129)
         );
  AOI22XL U60 ( .A0(n3), .A1(n127), .B0(n126), .B1(n131), .Y(n128) );
  OAI22XL U61 ( .A0(n3), .A1(n2), .B0(n4), .B1(n5), .Y(n124) );
  AOI222XL U62 ( .A0(n111), .A1(n126), .B0(n110), .B1(n14), .C0(n109), .C1(
        n108), .Y(n112) );
  OAI211XL U63 ( .A0(n107), .A1(n131), .B0(n2), .C0(addr[6]), .Y(n113) );
  OAI21XL U64 ( .A0(n1), .A1(addr[1]), .B0(n77), .Y(n81) );
  AOI221XL U65 ( .A0(n87), .A1(n14), .B0(n88), .B1(n126), .C0(n86), .Y(n90) );
  OAI211X1 U66 ( .A0(n85), .A1(n15), .B0(n84), .C0(n83), .Y(n86) );
  AOI222XL U67 ( .A0(n82), .A1(n14), .B0(n108), .B1(n107), .C0(n131), .C1(n79), 
        .Y(n85) );
  OAI21XL U68 ( .A0(n92), .A1(n13), .B0(addr[4]), .Y(n84) );
  AOI221XL U69 ( .A0(n126), .A1(n12), .B0(addr[3]), .B1(n127), .C0(n97), .Y(
        n98) );
  OAI22X1 U70 ( .A0(n18), .A1(n8), .B0(n5), .B1(n20), .Y(n97) );
  OAI211X1 U71 ( .A0(n78), .A1(n8), .B0(n119), .C0(n118), .Y(dout[3]) );
  AOI32XL U72 ( .A0(n126), .A1(n4), .A2(n103), .B0(n109), .B1(n110), .Y(n119)
         );
  AOI22XL U73 ( .A0(n117), .A1(n17), .B0(addr[5]), .B1(n116), .Y(n118) );
  AOI221XL U74 ( .A0(n122), .A1(n126), .B0(n96), .B1(n109), .C0(n10), .Y(n89)
         );
  AOI221XL U75 ( .A0(n131), .A1(n81), .B0(n95), .B1(n123), .C0(n80), .Y(n91)
         );
  NAND4X1 U76 ( .A(n102), .B(n114), .C(n101), .D(n100), .Y(dout[2]) );
  NAND3XL U77 ( .A(n3), .B(n125), .C(n103), .Y(n102) );
  AOI2BB2XL U78 ( .B0(addr[5]), .B1(n99), .A0N(addr[5]), .A1N(n98), .Y(n100)
         );
  OAI221X1 U79 ( .A0(n134), .A1(n17), .B0(n3), .B1(n133), .C0(n132), .Y(
        dout[4]) );
  AOI32XL U80 ( .A0(n131), .A1(n76), .A2(n1), .B0(n130), .B1(n17), .Y(n132) );
  AOI222XL U81 ( .A0(n12), .A1(n123), .B0(n122), .B1(addr[1]), .C0(n121), .C1(
        n19), .Y(n134) );
  CLKINVX3 U82 ( .A(n3), .Y(n7) );
  CLKINVX3 U83 ( .A(addr[3]), .Y(n14) );
endmodule


module sbox4_14 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126;

  OAI32X4 U12 ( .A0(n6), .A1(n2), .A2(addr[2]), .B0(n72), .B1(n108), .Y(n123)
         );
  OAI222X4 U20 ( .A0(addr[2]), .A1(n92), .B0(n106), .B1(n91), .C0(n90), .C1(
        n71), .Y(dout[2]) );
  OAI222X4 U33 ( .A0(addr[4]), .A1(n106), .B0(n16), .B1(n108), .C0(n2), .C1(
        n118), .Y(n83) );
  NAND2X2 U34 ( .A(addr[4]), .B(n2), .Y(n108) );
  NOR2X2 U43 ( .A(n8), .B(addr[4]), .Y(n113) );
  NOR2X2 U45 ( .A(n72), .B(n2), .Y(n111) );
  NAND2X2 U51 ( .A(n16), .B(n13), .Y(n118) );
  NOR2X2 U52 ( .A(n7), .B(addr[5]), .Y(n97) );
  NAND2X2 U53 ( .A(addr[6]), .B(addr[1]), .Y(n85) );
  NAND2X2 U54 ( .A(addr[1]), .B(n13), .Y(n116) );
  NOR2X2 U55 ( .A(n115), .B(n72), .Y(n121) );
  NAND2X2 U56 ( .A(n8), .B(n7), .Y(n115) );
  NAND2X2 U57 ( .A(addr[5]), .B(n7), .Y(n96) );
  NAND2X2 U58 ( .A(addr[6]), .B(n16), .Y(n106) );
  OAI222X1 U1 ( .A0(n6), .A1(n85), .B0(n97), .B1(n116), .C0(n7), .C1(n118), 
        .Y(n73) );
  CLKINVX1 U2 ( .A(n116), .Y(n12) );
  OAI31X4 U3 ( .A0(n118), .A1(n72), .A2(n7), .B0(n117), .Y(n119) );
  CLKINVX1 U4 ( .A(n8), .Y(n1) );
  CLKBUFX3 U5 ( .A(addr[3]), .Y(n2) );
  OAI221X1 U6 ( .A0(addr[2]), .A1(n80), .B0(n118), .B1(n105), .C0(n79), .Y(
        dout[1]) );
  AOI222XL U7 ( .A0(n7), .A1(n13), .B0(n113), .B1(n16), .C0(addr[1]), .C1(n8), 
        .Y(n114) );
  OAI222X1 U8 ( .A0(addr[1]), .A1(n84), .B0(n85), .B1(n74), .C0(n8), .C1(n107), 
        .Y(n75) );
  INVX4 U9 ( .A(addr[5]), .Y(n72) );
  OAI31X1 U10 ( .A0(n108), .A1(addr[5]), .A2(n14), .B0(n107), .Y(n109) );
  NAND2XL U11 ( .A(n1), .B(addr[5]), .Y(n84) );
  AOI211XL U13 ( .A0(n83), .A1(n72), .B0(n82), .C0(n5), .Y(n92) );
  NAND2XL U14 ( .A(n7), .B(n72), .Y(n74) );
  CLKINVX1 U15 ( .A(n118), .Y(n10) );
  CLKINVX1 U16 ( .A(n115), .Y(n4) );
  CLKINVX1 U17 ( .A(n112), .Y(n11) );
  OAI21X1 U18 ( .A0(n12), .A1(n14), .B0(n71), .Y(n112) );
  AOI22X1 U19 ( .A0(n15), .A1(n111), .B0(n14), .B1(n113), .Y(n93) );
  OAI211X1 U21 ( .A0(n16), .A1(n115), .B0(n93), .C0(n3), .Y(n94) );
  CLKINVX1 U22 ( .A(n85), .Y(n15) );
  NAND2X1 U23 ( .A(n97), .B(n8), .Y(n105) );
  NAND2X1 U24 ( .A(n113), .B(n10), .Y(n98) );
  NAND2X1 U25 ( .A(n12), .B(n97), .Y(n107) );
  NAND2X1 U26 ( .A(n118), .B(n85), .Y(n110) );
  OAI21XL U27 ( .A0(n4), .A1(n72), .B0(n108), .Y(n95) );
  CLKINVX1 U28 ( .A(n84), .Y(n9) );
  CLKINVX1 U29 ( .A(addr[2]), .Y(n71) );
  OAI31X1 U30 ( .A0(n7), .A1(addr[6]), .A2(n72), .B0(n87), .Y(n88) );
  OAI21XL U31 ( .A0(n113), .A1(n6), .B0(n15), .Y(n87) );
  OAI211X1 U32 ( .A0(n76), .A1(n7), .B0(n98), .C0(n3), .Y(n77) );
  AOI222XL U35 ( .A0(addr[5]), .A1(addr[6]), .B0(n111), .B1(addr[1]), .C0(n14), 
        .C1(n2), .Y(n76) );
  NAND3XL U36 ( .A(n15), .B(n8), .C(addr[4]), .Y(n117) );
  OAI22XL U37 ( .A0(n116), .A1(n115), .B0(n1), .B1(n112), .Y(n78) );
  CLKINVX3 U38 ( .A(addr[4]), .Y(n7) );
  OAI2BB2XL U39 ( .B0(n115), .B1(n106), .A0N(n72), .A1N(n86), .Y(n89) );
  OAI221XL U40 ( .A0(n116), .A1(addr[4]), .B0(n108), .B1(addr[1]), .C0(n117), 
        .Y(n86) );
  CLKINVX1 U41 ( .A(addr[6]), .Y(n13) );
  CLKINVX1 U42 ( .A(n81), .Y(n5) );
  OAI21XL U44 ( .A0(n96), .A1(n118), .B0(n93), .Y(n82) );
  NAND3X1 U46 ( .A(n101), .B(n100), .C(n99), .Y(n102) );
  AOI32X1 U47 ( .A0(n96), .A1(n8), .A2(n12), .B0(n15), .B1(n95), .Y(n101) );
  AOI2BB2XL U48 ( .B0(n16), .B1(n121), .A0N(n98), .A1N(addr[5]), .Y(n99) );
  OAI21XL U49 ( .A0(n97), .A1(n6), .B0(n14), .Y(n100) );
  AOI2BB2XL U50 ( .B0(n14), .B1(n123), .A0N(n122), .A1N(n71), .Y(n124) );
  AOI211XL U59 ( .A0(n14), .A1(n121), .B0(n120), .C0(n119), .Y(n122) );
  OAI22XL U60 ( .A0(n116), .A1(n115), .B0(addr[5]), .B1(n114), .Y(n120) );
  CLKINVX1 U61 ( .A(n75), .Y(n3) );
  AOI32XL U62 ( .A0(n12), .A1(n96), .A2(n1), .B0(addr[1]), .B1(n121), .Y(n81)
         );
  AOI222XL U63 ( .A0(n14), .A1(n6), .B0(n121), .B1(n116), .C0(n2), .C1(n73), 
        .Y(n80) );
  AOI22XL U64 ( .A0(n78), .A1(n72), .B0(addr[2]), .B1(n77), .Y(n79) );
  NAND2XL U65 ( .A(n111), .B(addr[4]), .Y(n91) );
  AOI211X1 U66 ( .A0(n9), .A1(n110), .B0(n89), .C0(n88), .Y(n90) );
  OAI211X1 U67 ( .A0(n106), .A1(n105), .B0(n104), .C0(n103), .Y(dout[3]) );
  AOI32X1 U68 ( .A0(n2), .A1(n6), .A2(n12), .B0(n94), .B1(n71), .Y(n104) );
  AOI22XL U69 ( .A0(addr[2]), .A1(n102), .B0(n10), .B1(n123), .Y(n103) );
  OAI211X1 U70 ( .A0(addr[2]), .A1(n126), .B0(n125), .C0(n124), .Y(dout[4]) );
  AOI32X1 U71 ( .A0(n15), .A1(n6), .A2(n2), .B0(n11), .B1(n9), .Y(n125) );
  AOI221XL U72 ( .A0(n10), .A1(n111), .B0(n4), .B1(n110), .C0(n109), .Y(n126)
         );
  CLKINVX3 U73 ( .A(n96), .Y(n6) );
  CLKINVX3 U74 ( .A(n2), .Y(n8) );
  CLKINVX3 U75 ( .A(n106), .Y(n14) );
  CLKINVX3 U76 ( .A(addr[1]), .Y(n16) );
endmodule


module sbox5_14 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121;

  OAI222X4 U18 ( .A0(addr[3]), .A1(n106), .B0(n14), .B1(n90), .C0(n5), .C1(n70), .Y(n93) );
  OAI22X2 U40 ( .A0(addr[5]), .A1(n106), .B0(n68), .B1(n114), .Y(n116) );
  NOR2X2 U41 ( .A(n3), .B(addr[3]), .Y(n102) );
  NAND2X2 U45 ( .A(addr[6]), .B(n70), .Y(n114) );
  NAND2X2 U50 ( .A(n70), .B(n14), .Y(n110) );
  NAND2X2 U52 ( .A(addr[1]), .B(n14), .Y(n113) );
  NAND2X2 U54 ( .A(addr[1]), .B(addr[6]), .Y(n106) );
  NAND2X2 U55 ( .A(addr[3]), .B(n5), .Y(n121) );
  CLKINVX1 U1 ( .A(addr[5]), .Y(n1) );
  AOI221XL U2 ( .A0(n93), .A1(n1), .B0(n15), .B1(n7), .C0(n92), .Y(n105) );
  INVX3 U3 ( .A(addr[5]), .Y(n68) );
  OAI221X4 U4 ( .A0(n111), .A1(n110), .B0(n121), .B1(n114), .C0(n109), .Y(n112) );
  OAI221X4 U5 ( .A0(n5), .A1(n114), .B0(n68), .B1(n113), .C0(n120), .Y(n115)
         );
  OAI221X4 U6 ( .A0(n107), .A1(n121), .B0(n111), .B1(n113), .C0(n85), .Y(n86)
         );
  OAI31X1 U7 ( .A0(n9), .A1(addr[5]), .A2(addr[1]), .B0(n81), .Y(n73) );
  OAI32X1 U8 ( .A0(n114), .A1(addr[5]), .A2(n3), .B0(n4), .B1(n107), .Y(n79)
         );
  AOI32XL U9 ( .A0(n7), .A1(n98), .A2(n13), .B0(n2), .B1(n73), .Y(n77) );
  CLKBUFX3 U10 ( .A(addr[4]), .Y(n2) );
  CLKINVX1 U11 ( .A(n81), .Y(n6) );
  NAND2X1 U12 ( .A(n16), .B(n7), .Y(n81) );
  CLKINVX1 U13 ( .A(n110), .Y(n11) );
  CLKXOR2X2 U14 ( .A(n9), .B(n68), .Y(n94) );
  AOI2BB1X1 U15 ( .A0N(n5), .A1N(n1), .B0(n7), .Y(n111) );
  NOR2X1 U16 ( .A(n121), .B(n68), .Y(n91) );
  NOR2BX1 U17 ( .AN(n116), .B(n90), .Y(n83) );
  NAND2X1 U19 ( .A(n11), .B(n68), .Y(n120) );
  CLKINVX1 U20 ( .A(n113), .Y(n13) );
  NAND2X1 U21 ( .A(n13), .B(n68), .Y(n107) );
  CLKINVX1 U22 ( .A(n121), .Y(n4) );
  OAI31X1 U23 ( .A0(n69), .A1(n7), .A2(n113), .B0(n99), .Y(n72) );
  CLKINVX1 U24 ( .A(n106), .Y(n15) );
  OAI2BB2XL U25 ( .B0(n1), .B1(n113), .A0N(n98), .A1N(n16), .Y(n101) );
  CLKINVX1 U26 ( .A(n114), .Y(n16) );
  CLKINVX1 U27 ( .A(n90), .Y(n8) );
  CLKINVX1 U28 ( .A(addr[1]), .Y(n70) );
  CLKINVX1 U29 ( .A(addr[3]), .Y(n9) );
  CLKINVX1 U30 ( .A(addr[6]), .Y(n14) );
  AOI211X1 U31 ( .A0(n91), .A1(addr[1]), .B0(n80), .C0(n79), .Y(n89) );
  OAI2BB2XL U32 ( .B0(n111), .B1(n106), .A0N(n94), .A1N(n11), .Y(n80) );
  AOI211X1 U33 ( .A0(n102), .A1(n84), .B0(n83), .C0(n82), .Y(n85) );
  OAI21XL U34 ( .A0(n14), .A1(n1), .B0(n106), .Y(n84) );
  NOR3XL U35 ( .A(n94), .B(n3), .C(n110), .Y(n82) );
  AOI222XL U36 ( .A0(n15), .A1(n8), .B0(addr[5]), .B1(n108), .C0(n12), .C1(n5), 
        .Y(n109) );
  CLKINVX1 U37 ( .A(n107), .Y(n12) );
  OAI21XL U38 ( .A0(addr[6]), .A1(addr[3]), .B0(n106), .Y(n108) );
  NAND2X1 U39 ( .A(addr[3]), .B(n3), .Y(n90) );
  NAND2X1 U42 ( .A(n2), .B(addr[5]), .Y(n98) );
  NAND2X1 U43 ( .A(n3), .B(n9), .Y(n97) );
  OAI21XL U44 ( .A0(addr[1]), .A1(n97), .B0(n96), .Y(n103) );
  AOI33XL U46 ( .A0(n3), .A1(n95), .A2(addr[5]), .B0(n94), .B1(n5), .B2(
        addr[1]), .Y(n96) );
  OAI21XL U47 ( .A0(n70), .A1(n9), .B0(n114), .Y(n95) );
  OAI21XL U48 ( .A0(addr[6]), .A1(n121), .B0(n99), .Y(n100) );
  NAND2X1 U49 ( .A(n71), .B(n11), .Y(n99) );
  XOR2X1 U51 ( .A(n69), .B(n3), .Y(n71) );
  AOI2BB2XL U53 ( .B0(n102), .B1(n116), .A0N(n2), .A1N(n75), .Y(n76) );
  AOI211X1 U56 ( .A0(n10), .A1(n3), .B0(n74), .C0(n83), .Y(n75) );
  AO22XL U57 ( .A0(n13), .A1(n4), .B0(addr[6]), .B1(n102), .Y(n74) );
  CLKINVX1 U58 ( .A(n120), .Y(n10) );
  CLKINVX1 U59 ( .A(n2), .Y(n69) );
  AO22XL U60 ( .A0(n13), .A1(n8), .B0(addr[6]), .B1(n91), .Y(n92) );
  AOI222XL U61 ( .A0(n116), .A1(n5), .B0(addr[3]), .B1(n115), .C0(n13), .C1(n7), .Y(n117) );
  OAI221X1 U62 ( .A0(n2), .A1(n105), .B0(n110), .B1(n121), .C0(n104), .Y(
        dout[3]) );
  AOI222XL U63 ( .A0(n2), .A1(n103), .B0(n102), .B1(n101), .C0(n100), .C1(n1), 
        .Y(n104) );
  OAI211X1 U64 ( .A0(n2), .A1(n89), .B0(n88), .C0(n87), .Y(dout[2]) );
  AOI33XL U65 ( .A0(n4), .A1(n98), .A2(n16), .B0(n3), .B1(n94), .B2(n11), .Y(
        n88) );
  AOI222XL U66 ( .A0(n6), .A1(n68), .B0(n2), .B1(n86), .C0(n91), .C1(n15), .Y(
        n87) );
  OAI211X1 U67 ( .A0(n78), .A1(n68), .B0(n77), .C0(n76), .Y(dout[1]) );
  AOI221XL U68 ( .A0(n4), .A1(addr[1]), .B0(n15), .B1(n7), .C0(n72), .Y(n78)
         );
  OAI211X1 U69 ( .A0(n121), .A1(n120), .B0(n119), .C0(n118), .Y(dout[4]) );
  AOI32XL U70 ( .A0(n7), .A1(n114), .A2(addr[5]), .B0(n2), .B1(n112), .Y(n119)
         );
  AOI2BB2X1 U71 ( .B0(n6), .B1(n68), .A0N(n2), .A1N(n117), .Y(n118) );
  BUFX4 U72 ( .A(addr[2]), .Y(n3) );
  CLKINVX3 U73 ( .A(n3), .Y(n5) );
  CLKINVX3 U74 ( .A(n97), .Y(n7) );
endmodule


module sbox6_14 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147;

  NAND2X2 U39 ( .A(n138), .B(addr[3]), .Y(n147) );
  NOR2X2 U47 ( .A(n15), .B(n13), .Y(n138) );
  NOR2X2 U50 ( .A(n81), .B(n4), .Y(n119) );
  NOR2X2 U58 ( .A(n84), .B(n81), .Y(n125) );
  NAND2X2 U61 ( .A(n97), .B(n103), .Y(n112) );
  NOR2X2 U62 ( .A(n11), .B(addr[1]), .Y(n103) );
  NOR2X2 U63 ( .A(n84), .B(addr[3]), .Y(n97) );
  NAND2X2 U64 ( .A(n117), .B(n131), .Y(n140) );
  NOR2X2 U65 ( .A(n5), .B(addr[3]), .Y(n131) );
  NOR2X2 U66 ( .A(n83), .B(addr[6]), .Y(n117) );
  NOR2X1 U1 ( .A(n15), .B(addr[3]), .Y(n102) );
  OAI222X1 U2 ( .A0(n91), .A1(n85), .B0(n3), .B1(n82), .C0(addr[5]), .C1(n17), 
        .Y(n92) );
  CLKINVX1 U3 ( .A(addr[3]), .Y(n1) );
  INVX3 U4 ( .A(addr[3]), .Y(n81) );
  CLKINVX1 U5 ( .A(n84), .Y(n2) );
  INVX4 U6 ( .A(n4), .Y(n84) );
  CLKBUFX3 U7 ( .A(addr[4]), .Y(n4) );
  OAI221X1 U8 ( .A0(n11), .A1(n18), .B0(n81), .B1(n8), .C0(n86), .Y(n90) );
  CLKINVX1 U9 ( .A(n15), .Y(n3) );
  BUFX4 U10 ( .A(addr[2]), .Y(n5) );
  NOR2X4 U11 ( .A(addr[1]), .B(addr[6]), .Y(n130) );
  OAI22X1 U12 ( .A0(n81), .A1(n11), .B0(addr[1]), .B1(n17), .Y(n142) );
  OAI221X4 U13 ( .A0(n123), .A1(n10), .B0(n13), .B1(n85), .C0(n7), .Y(n124) );
  NOR2X4 U14 ( .A(n5), .B(addr[5]), .Y(n143) );
  INVX1 U15 ( .A(n130), .Y(n14) );
  CLKINVX1 U16 ( .A(n125), .Y(n18) );
  NAND2X1 U17 ( .A(n14), .B(n8), .Y(n105) );
  INVXL U18 ( .A(n121), .Y(n16) );
  CLKINVX1 U19 ( .A(n138), .Y(n12) );
  AOI211X1 U20 ( .A0(n85), .A1(n81), .B0(n131), .C0(n143), .Y(n121) );
  CLKINVX1 U21 ( .A(n117), .Y(n13) );
  CLKINVX1 U22 ( .A(n119), .Y(n17) );
  NOR2X1 U23 ( .A(n8), .B(n123), .Y(n144) );
  NOR2X1 U24 ( .A(n83), .B(n11), .Y(n96) );
  CLKINVX1 U25 ( .A(n103), .Y(n10) );
  OAI211X1 U26 ( .A0(n14), .A1(n18), .B0(n104), .C0(n112), .Y(n108) );
  OAI21XL U27 ( .A0(n103), .A1(n117), .B0(n102), .Y(n104) );
  OAI21XL U28 ( .A0(n132), .A1(n11), .B0(n1), .Y(n86) );
  AOI21X1 U29 ( .A0(n84), .A1(n102), .B0(n125), .Y(n91) );
  OAI2BB2XL U30 ( .B0(n143), .B1(n14), .A0N(n143), .A1N(n117), .Y(n118) );
  CLKINVX1 U31 ( .A(n122), .Y(n7) );
  CLKINVX1 U32 ( .A(n126), .Y(n9) );
  CLKINVX1 U33 ( .A(n97), .Y(n82) );
  NAND2BX1 U34 ( .AN(n144), .B(n137), .Y(n107) );
  CLKINVX1 U35 ( .A(addr[1]), .Y(n83) );
  NOR2X1 U36 ( .A(n8), .B(n3), .Y(n122) );
  NOR2X1 U37 ( .A(addr[1]), .B(n2), .Y(n132) );
  OAI22X1 U38 ( .A0(n17), .A1(n13), .B0(n5), .B1(n9), .Y(n88) );
  NAND2X1 U40 ( .A(n5), .B(n85), .Y(n123) );
  NAND4X1 U41 ( .A(n147), .B(n140), .C(n100), .D(n99), .Y(n101) );
  AOI222XL U42 ( .A0(n98), .A1(n15), .B0(n102), .B1(n130), .C0(n97), .C1(n105), 
        .Y(n99) );
  NAND3X1 U43 ( .A(n5), .B(n17), .C(n96), .Y(n100) );
  OAI221X1 U44 ( .A0(n81), .A1(n10), .B0(n17), .B1(n11), .C0(n9), .Y(n98) );
  AOI22X1 U45 ( .A0(n4), .A1(n115), .B0(addr[5]), .B1(n114), .Y(n129) );
  OAI21XL U46 ( .A0(n121), .A1(n14), .B0(n147), .Y(n115) );
  OAI21XL U48 ( .A0(n113), .A1(n15), .B0(n112), .Y(n114) );
  AOI221XL U49 ( .A0(n119), .A1(n83), .B0(n130), .B1(addr[3]), .C0(n111), .Y(
        n113) );
  OAI22XL U51 ( .A0(n13), .A1(n84), .B0(addr[3]), .B1(n8), .Y(n111) );
  AOI211X1 U52 ( .A0(n4), .A1(n135), .B0(n134), .C0(n133), .Y(n136) );
  OA21XL U53 ( .A0(n1), .A1(n3), .B0(n132), .Y(n133) );
  OAI2BB2XL U54 ( .B0(n2), .B1(n7), .A0N(n131), .A1N(n130), .Y(n134) );
  OAI22X1 U55 ( .A0(n5), .A1(n13), .B0(n15), .B1(n8), .Y(n135) );
  CLKINVX3 U56 ( .A(addr[5]), .Y(n85) );
  AOI2BB2X1 U57 ( .B0(n5), .B1(n130), .A0N(n3), .A1N(n10), .Y(n137) );
  NOR2X1 U59 ( .A(n10), .B(n2), .Y(n126) );
  AOI2BB2XL U60 ( .B0(n143), .B1(n90), .A0N(n89), .A1N(n85), .Y(n94) );
  AOI211X1 U67 ( .A0(n122), .A1(n4), .B0(n88), .C0(n87), .Y(n89) );
  OAI32X1 U68 ( .A0(n10), .A1(n81), .A2(n15), .B0(n12), .B1(n82), .Y(n87) );
  NAND3X1 U69 ( .A(n147), .B(n140), .C(n139), .Y(n141) );
  AOI32X1 U70 ( .A0(n5), .A1(n83), .A2(n4), .B0(n138), .B1(n84), .Y(n139) );
  AO22XL U71 ( .A0(n143), .A1(n2), .B0(n116), .B1(n84), .Y(n120) );
  OAI21XL U72 ( .A0(n3), .A1(n85), .B0(n123), .Y(n116) );
  CLKINVX1 U73 ( .A(n106), .Y(n6) );
  AOI32XL U74 ( .A0(n105), .A1(n84), .A2(n1), .B0(addr[1]), .B1(n125), .Y(n106) );
  OAI211X1 U75 ( .A0(n84), .A1(n140), .B0(n110), .C0(n109), .Y(dout[2]) );
  AOI222XL U76 ( .A0(n108), .A1(n85), .B0(n143), .B1(n6), .C0(n119), .C1(n107), 
        .Y(n109) );
  AOI2BB2XL U77 ( .B0(addr[5]), .B1(n101), .A0N(n15), .A1N(n112), .Y(n110) );
  OAI211X1 U78 ( .A0(n2), .A1(n147), .B0(n146), .C0(n145), .Y(dout[4]) );
  AOI222XL U79 ( .A0(n144), .A1(n81), .B0(n143), .B1(n142), .C0(n141), .C1(n85), .Y(n145) );
  OA22X1 U80 ( .A0(n18), .A1(n137), .B0(n136), .B1(n85), .Y(n146) );
  NAND3X1 U81 ( .A(n129), .B(n128), .C(n127), .Y(dout[3]) );
  AOI32XL U82 ( .A0(n120), .A1(n81), .A2(addr[1]), .B0(n119), .B1(n118), .Y(
        n128) );
  AOI222XL U83 ( .A0(n144), .A1(n84), .B0(n126), .B1(n16), .C0(n125), .C1(n124), .Y(n127) );
  NAND3BX1 U84 ( .AN(n95), .B(n94), .C(n93), .Y(dout[1]) );
  OAI222X1 U85 ( .A0(n140), .A1(n4), .B0(n112), .B1(n15), .C0(n8), .C1(n91), 
        .Y(n95) );
  AOI32XL U86 ( .A0(addr[1]), .A1(n85), .A2(n125), .B0(n130), .B1(n92), .Y(n93) );
  CLKINVX3 U87 ( .A(n96), .Y(n8) );
  CLKINVX3 U88 ( .A(addr[6]), .Y(n11) );
  CLKINVX3 U89 ( .A(n5), .Y(n15) );
endmodule


module sbox7_14 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148;

  OAI222X4 U19 ( .A0(n20), .A1(n129), .B0(n4), .B1(n13), .C0(addr[1]), .C1(n12), .Y(n122) );
  OAI33X4 U33 ( .A0(addr[1]), .A1(n4), .A2(n5), .B0(n18), .B1(n21), .B2(n6), 
        .Y(n97) );
  NOR2X2 U44 ( .A(n10), .B(n4), .Y(n116) );
  NOR2X2 U48 ( .A(addr[1]), .B(addr[6]), .Y(n136) );
  NOR2X2 U51 ( .A(n87), .B(n10), .Y(n125) );
  NOR2X2 U52 ( .A(n18), .B(addr[3]), .Y(n131) );
  NOR2X2 U58 ( .A(n93), .B(n124), .Y(n142) );
  NOR2X2 U60 ( .A(n19), .B(addr[1]), .Y(n93) );
  NOR2X2 U62 ( .A(n84), .B(n3), .Y(n137) );
  NOR2X2 U65 ( .A(n19), .B(n86), .Y(n140) );
  NAND2X1 U1 ( .A(n3), .B(n4), .Y(n119) );
  CLKBUFX3 U2 ( .A(addr[4]), .Y(n4) );
  CLKINVX1 U3 ( .A(n84), .Y(n1) );
  CLKINVX1 U4 ( .A(n21), .Y(n2) );
  CLKBUFX3 U5 ( .A(addr[2]), .Y(n5) );
  OAI31X1 U6 ( .A0(n10), .A1(n84), .A2(n86), .B0(n117), .Y(n121) );
  NOR2X4 U7 ( .A(n86), .B(addr[6]), .Y(n124) );
  OAI22X1 U8 ( .A0(addr[1]), .A1(n12), .B0(n5), .B1(n113), .Y(n100) );
  OAI22X1 U9 ( .A0(n4), .A1(n87), .B0(addr[3]), .B1(n83), .Y(n103) );
  AOI211XL U10 ( .A0(n5), .A1(n17), .B0(n131), .C0(n130), .Y(n132) );
  NOR3XL U11 ( .A(n20), .B(addr[3]), .C(n2), .Y(n130) );
  OAI21XL U12 ( .A0(n3), .A1(n1), .B0(n119), .Y(n89) );
  BUFX4 U13 ( .A(addr[5]), .Y(n3) );
  AOI221XL U14 ( .A0(n140), .A1(n89), .B0(n109), .B1(n17), .C0(n88), .Y(n96)
         );
  CLKINVX1 U15 ( .A(n140), .Y(n18) );
  OAI2BB2XL U16 ( .B0(n142), .B1(n83), .A0N(n141), .A1N(n140), .Y(n143) );
  CLKINVX1 U17 ( .A(n125), .Y(n8) );
  CLKINVX1 U18 ( .A(n142), .Y(n17) );
  NAND2X1 U20 ( .A(n8), .B(n14), .Y(n105) );
  CLKINVX1 U21 ( .A(n123), .Y(n11) );
  CLKINVX1 U22 ( .A(n109), .Y(n9) );
  NAND2X1 U23 ( .A(n124), .B(n10), .Y(n113) );
  CLKINVX1 U24 ( .A(n137), .Y(n83) );
  NOR2X1 U25 ( .A(n83), .B(n10), .Y(n109) );
  CLKINVX1 U26 ( .A(n136), .Y(n20) );
  OAI22XL U27 ( .A0(n137), .A1(n13), .B0(n86), .B1(n9), .Y(n146) );
  OAI21X1 U28 ( .A0(n84), .A1(n8), .B0(n129), .Y(n141) );
  NAND2X1 U29 ( .A(n116), .B(n87), .Y(n129) );
  CLKINVX1 U30 ( .A(n93), .Y(n16) );
  OAI21XL U31 ( .A0(n119), .A1(n16), .B0(n118), .Y(n120) );
  OAI21XL U32 ( .A0(n125), .A1(n137), .B0(n124), .Y(n118) );
  NOR2X1 U34 ( .A(n87), .B(n12), .Y(n123) );
  CLKINVX1 U35 ( .A(n145), .Y(n12) );
  OAI22XL U36 ( .A0(n137), .A1(n113), .B0(n19), .B1(n11), .Y(n88) );
  CLKINVX1 U37 ( .A(n116), .Y(n6) );
  CLKINVX1 U38 ( .A(n131), .Y(n13) );
  CLKINVX1 U39 ( .A(n134), .Y(n14) );
  NOR2XL U40 ( .A(n125), .B(n84), .Y(n110) );
  CLKINVX1 U41 ( .A(n119), .Y(n85) );
  CLKINVX1 U42 ( .A(n103), .Y(n15) );
  OA21XL U43 ( .A0(n7), .A1(n16), .B0(n117), .Y(n102) );
  CLKINVX1 U45 ( .A(n105), .Y(n7) );
  OAI2BB1XL U46 ( .A0N(n103), .A1N(n124), .B0(n102), .Y(n104) );
  OAI22X1 U47 ( .A0(n87), .A1(n6), .B0(n4), .B1(n14), .Y(n112) );
  NOR4X1 U49 ( .A(n4), .B(addr[3]), .C(n86), .D(n21), .Y(n99) );
  XNOR2X1 U50 ( .A(addr[6]), .B(n5), .Y(n101) );
  AOI211X1 U53 ( .A0(n116), .A1(addr[6]), .B0(n115), .C0(n114), .Y(n128) );
  OAI222X1 U54 ( .A0(n111), .A1(n18), .B0(n110), .B1(n16), .C0(n20), .C1(n9), 
        .Y(n115) );
  OAI2BB2XL U55 ( .B0(n85), .B1(n113), .A0N(n86), .A1N(n112), .Y(n114) );
  OA21XL U56 ( .A0(n10), .A1(n3), .B0(n11), .Y(n111) );
  NAND2X1 U57 ( .A(n5), .B(n136), .Y(n133) );
  CLKINVX1 U59 ( .A(addr[6]), .Y(n19) );
  AOI211X1 U61 ( .A0(n131), .A1(n3), .B0(n92), .C0(n91), .Y(n95) );
  OAI221X1 U63 ( .A0(n86), .A1(n12), .B0(n18), .B1(n83), .C0(n102), .Y(n92) );
  OAI31X1 U64 ( .A0(n10), .A1(n84), .A2(n20), .B0(n90), .Y(n91) );
  AO21XL U66 ( .A0(n119), .A1(n129), .B0(addr[6]), .Y(n90) );
  NOR2X1 U67 ( .A(n84), .B(addr[3]), .Y(n145) );
  AOI21XL U68 ( .A0(addr[3]), .A1(n98), .B0(n97), .Y(n108) );
  OAI2BB1XL U69 ( .A0N(n21), .A1N(n124), .B0(n133), .Y(n98) );
  NAND3X1 U70 ( .A(n136), .B(n10), .C(n3), .Y(n117) );
  NOR2X1 U71 ( .A(addr[3]), .B(n3), .Y(n134) );
  OAI21X1 U72 ( .A0(n5), .A1(n142), .B0(n133), .Y(n138) );
  OAI22XL U73 ( .A0(n142), .A1(n6), .B0(n1), .B1(n132), .Y(n135) );
  AO21X1 U74 ( .A0(n139), .A1(n87), .B0(n138), .Y(n144) );
  OAI21XL U75 ( .A0(n2), .A1(n86), .B0(n16), .Y(n139) );
  OAI221X1 U76 ( .A0(n96), .A1(n21), .B0(n5), .B1(n95), .C0(n94), .Y(dout[1])
         );
  AOI2BB2X1 U77 ( .B0(n93), .B1(n112), .A0N(n133), .A1N(n15), .Y(n94) );
  OAI211X1 U78 ( .A0(n128), .A1(n21), .B0(n127), .C0(n126), .Y(dout[3]) );
  AOI32XL U79 ( .A0(n125), .A1(n1), .A2(n124), .B0(n123), .B1(n136), .Y(n126)
         );
  OAI31X1 U80 ( .A0(n122), .A1(n121), .A2(n120), .B0(n21), .Y(n127) );
  OAI221X1 U81 ( .A0(n3), .A1(n108), .B0(n107), .B1(n87), .C0(n106), .Y(
        dout[2]) );
  AOI32XL U82 ( .A0(n105), .A1(n21), .A2(n140), .B0(n2), .B1(n104), .Y(n106)
         );
  AOI211X1 U83 ( .A0(n101), .A1(n4), .B0(n100), .C0(n99), .Y(n107) );
  NAND2X1 U84 ( .A(n148), .B(n147), .Y(dout[4]) );
  AOI222XL U85 ( .A0(n136), .A1(n141), .B0(n3), .B1(n135), .C0(n134), .C1(n138), .Y(n148) );
  AOI222XL U86 ( .A0(n5), .A1(n146), .B0(n145), .B1(n144), .C0(n143), .C1(n21), 
        .Y(n147) );
  CLKINVX3 U87 ( .A(addr[3]), .Y(n10) );
  CLKINVX3 U88 ( .A(n5), .Y(n21) );
  CLKINVX3 U89 ( .A(n4), .Y(n84) );
  CLKINVX3 U90 ( .A(addr[1]), .Y(n86) );
  CLKINVX3 U91 ( .A(n3), .Y(n87) );
endmodule


module sbox8_14 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132;

  NAND2X2 U41 ( .A(addr[6]), .B(n10), .Y(n131) );
  NAND2X2 U48 ( .A(addr[4]), .B(n13), .Y(n123) );
  NAND2X2 U49 ( .A(n2), .B(n74), .Y(n87) );
  NAND2X2 U50 ( .A(addr[1]), .B(n6), .Y(n124) );
  NAND2X2 U54 ( .A(addr[2]), .B(n15), .Y(n116) );
  NAND2X2 U60 ( .A(addr[6]), .B(addr[1]), .Y(n105) );
  NAND2X2 U61 ( .A(n10), .B(n6), .Y(n108) );
  OAI32X1 U1 ( .A0(n6), .A1(addr[4]), .A2(n92), .B0(n115), .B1(n108), .Y(n96)
         );
  OAI31X1 U2 ( .A0(n123), .A1(addr[6]), .A2(n116), .B0(n109), .Y(n110) );
  AOI222X1 U3 ( .A0(n88), .A1(addr[2]), .B0(n74), .B1(n16), .C0(n75), .C1(n92), 
        .Y(n114) );
  OAI222X1 U4 ( .A0(addr[2]), .A1(n126), .B0(n13), .B1(n125), .C0(n124), .C1(
        n123), .Y(n127) );
  OAI221X1 U5 ( .A0(n105), .A1(n87), .B0(addr[4]), .B1(n108), .C0(n86), .Y(n90) );
  NAND2X4 U6 ( .A(addr[4]), .B(n2), .Y(n115) );
  AOI32XL U7 ( .A0(n4), .A1(n14), .A2(n2), .B0(n5), .B1(n117), .Y(n130) );
  OA21XL U8 ( .A0(n75), .A1(n15), .B0(n121), .Y(n78) );
  INVXL U9 ( .A(n119), .Y(n3) );
  INVX3 U10 ( .A(n2), .Y(n13) );
  BUFX4 U11 ( .A(addr[3]), .Y(n2) );
  CLKBUFX3 U12 ( .A(addr[5]), .Y(n1) );
  CLKINVX1 U13 ( .A(n108), .Y(n5) );
  CLKINVX1 U14 ( .A(n107), .Y(n11) );
  CLKINVX1 U15 ( .A(n93), .Y(n12) );
  NAND2X1 U16 ( .A(n13), .B(n74), .Y(n93) );
  NAND2X1 U17 ( .A(n75), .B(n15), .Y(n121) );
  OAI21XL U18 ( .A0(n115), .A1(n15), .B0(n107), .Y(n77) );
  OAI21X1 U19 ( .A0(n74), .A1(n15), .B0(n123), .Y(n88) );
  OAI31XL U20 ( .A0(n115), .A1(n10), .A2(n116), .B0(n118), .Y(n94) );
  CLKINVX1 U21 ( .A(n131), .Y(n9) );
  NAND2X1 U22 ( .A(n14), .B(n13), .Y(n107) );
  OAI22XL U23 ( .A0(n116), .A1(n123), .B0(n14), .B1(n115), .Y(n117) );
  OAI22XL U24 ( .A0(n123), .A1(n108), .B0(n131), .B1(n93), .Y(n95) );
  OAI2BB2XL U25 ( .B0(n115), .B1(n131), .A0N(n88), .A1N(n8), .Y(n89) );
  AOI211XL U26 ( .A0(n108), .A1(n105), .B0(n74), .C0(n121), .Y(n85) );
  CLKINVX1 U27 ( .A(n124), .Y(n4) );
  OAI22XL U28 ( .A0(n14), .A1(n123), .B0(n78), .B1(n87), .Y(n81) );
  NAND2BX2 U29 ( .AN(n78), .B(n13), .Y(n120) );
  NAND2XL U30 ( .A(n115), .B(n93), .Y(n104) );
  OAI2BB2XL U31 ( .B0(n106), .B1(n105), .A0N(n104), .A1N(n4), .Y(n111) );
  NOR2BXL U32 ( .AN(n123), .B(n103), .Y(n106) );
  NAND3X1 U33 ( .A(n104), .B(n10), .C(n14), .Y(n84) );
  AO21X1 U34 ( .A0(n14), .A1(n8), .B0(n101), .Y(n102) );
  OAI33X1 U35 ( .A0(n6), .A1(n13), .A2(n100), .B0(n75), .B1(n103), .B2(n124), 
        .Y(n101) );
  OA22XL U36 ( .A0(n107), .A1(n131), .B0(n120), .B1(n124), .Y(n98) );
  CLKINVX1 U37 ( .A(n125), .Y(n7) );
  OAI21XL U38 ( .A0(n4), .A1(n9), .B0(addr[4]), .Y(n86) );
  NAND2X1 U39 ( .A(n1), .B(n75), .Y(n100) );
  OAI221X1 U40 ( .A0(n124), .A1(n121), .B0(addr[1]), .B1(n120), .C0(n3), .Y(
        n128) );
  OAI31XL U42 ( .A0(n75), .A1(n10), .A2(n13), .B0(n118), .Y(n119) );
  NAND2X1 U43 ( .A(n8), .B(addr[2]), .Y(n125) );
  NAND4XL U44 ( .A(n9), .B(n1), .C(n2), .D(addr[2]), .Y(n109) );
  NAND3X1 U45 ( .A(n14), .B(n6), .C(n2), .Y(n118) );
  OAI21XL U46 ( .A0(n1), .A1(n87), .B0(n114), .Y(n76) );
  OAI22XL U47 ( .A0(n108), .A1(n120), .B0(n79), .B1(n100), .Y(n80) );
  AOI221XL U51 ( .A0(n9), .A1(n13), .B0(n8), .B1(n2), .C0(n91), .Y(n79) );
  NOR2X1 U52 ( .A(n1), .B(n2), .Y(n103) );
  NOR2X1 U53 ( .A(n87), .B(addr[6]), .Y(n91) );
  NOR2X1 U55 ( .A(n13), .B(n1), .Y(n92) );
  CLKINVX1 U56 ( .A(n100), .Y(n16) );
  OA21XL U57 ( .A0(n1), .A1(n115), .B0(n120), .Y(n132) );
  AOI221XL U58 ( .A0(n5), .A1(n2), .B0(n8), .B1(addr[4]), .C0(n122), .Y(n126)
         );
  OAI22XL U59 ( .A0(n2), .A1(n10), .B0(addr[4]), .B1(n131), .Y(n122) );
  OAI211X1 U62 ( .A0(addr[2]), .A1(n99), .B0(n98), .C0(n97), .Y(dout[2]) );
  AOI221XL U63 ( .A0(addr[2]), .A1(n96), .B0(n1), .B1(n95), .C0(n94), .Y(n97)
         );
  AOI221XL U64 ( .A0(n91), .A1(n1), .B0(n90), .B1(n15), .C0(n89), .Y(n99) );
  OAI211X1 U65 ( .A0(n132), .A1(n131), .B0(n130), .C0(n129), .Y(dout[4]) );
  AOI222XL U66 ( .A0(n128), .A1(n74), .B0(n1), .B1(n127), .C0(n11), .C1(n8), 
        .Y(n129) );
  OAI211X1 U67 ( .A0(addr[1]), .A1(n114), .B0(n113), .C0(n112), .Y(dout[3]) );
  AOI221XL U68 ( .A0(n111), .A1(n75), .B0(n11), .B1(n5), .C0(n110), .Y(n112)
         );
  AOI2BB2XL U69 ( .B0(n102), .B1(n74), .A0N(n115), .A1N(n125), .Y(n113) );
  NAND4BX1 U70 ( .AN(n85), .B(n84), .C(n83), .D(n82), .Y(dout[1]) );
  AOI221XL U71 ( .A0(n9), .A1(n81), .B0(n12), .B1(n7), .C0(n80), .Y(n82) );
  AOI22X1 U72 ( .A0(n8), .A1(n77), .B0(n4), .B1(n76), .Y(n83) );
  CLKINVX3 U73 ( .A(addr[6]), .Y(n6) );
  CLKINVX3 U74 ( .A(n105), .Y(n8) );
  CLKINVX3 U75 ( .A(addr[1]), .Y(n10) );
  CLKINVX3 U76 ( .A(n116), .Y(n14) );
  CLKINVX3 U77 ( .A(n1), .Y(n15) );
  CLKINVX3 U78 ( .A(addr[4]), .Y(n74) );
  CLKINVX3 U79 ( .A(addr[2]), .Y(n75) );
endmodule


module crp_14 ( P, R, K_sub );
  output [1:32] P;
  input [1:32] R;
  input [1:48] K_sub;
  wire   n1;
  wire   [1:48] X;

  sbox1_14 u0 ( .addr(X[1:6]), .dout({P[9], P[17], P[23], P[31]}) );
  sbox2_14 u1 ( .addr({X[7], n1, X[9:12]}), .dout({P[13], P[28], P[2], P[18]})
         );
  sbox3_14 u2 ( .addr(X[13:18]), .dout({P[24], P[16], P[30], P[6]}) );
  sbox4_14 u3 ( .addr(X[19:24]), .dout({P[26], P[20], P[10], P[1]}) );
  sbox5_14 u4 ( .addr(X[25:30]), .dout({P[8], P[14], P[25], P[3]}) );
  sbox6_14 u5 ( .addr(X[31:36]), .dout({P[4], P[29], P[11], P[19]}) );
  sbox7_14 u6 ( .addr(X[37:42]), .dout({P[32], P[12], P[22], P[7]}) );
  sbox8_14 u7 ( .addr(X[43:48]), .dout({P[5], P[27], P[15], P[21]}) );
  XOR2X1 U1 ( .A(R[1]), .B(K_sub[2]), .Y(X[2]) );
  CLKXOR2X4 U2 ( .A(R[10]), .B(K_sub[15]), .Y(X[15]) );
  CLKXOR2X4 U3 ( .A(R[8]), .B(K_sub[11]), .Y(X[11]) );
  CLKXOR2X4 U4 ( .A(R[29]), .B(K_sub[42]), .Y(X[42]) );
  CLKXOR2X4 U5 ( .A(R[5]), .B(K_sub[6]), .Y(X[6]) );
  CLKXOR2X4 U6 ( .A(R[20]), .B(K_sub[31]), .Y(X[31]) );
  CLKXOR2X4 U7 ( .A(R[16]), .B(K_sub[25]), .Y(X[25]) );
  CLKXOR2X4 U8 ( .A(R[29]), .B(K_sub[44]), .Y(X[44]) );
  CLKXOR2X4 U9 ( .A(R[12]), .B(K_sub[19]), .Y(X[19]) );
  XNOR2X1 U10 ( .A(R[5]), .B(K_sub[8]), .Y(X[8]) );
  INVX3 U11 ( .A(X[8]), .Y(n1) );
  CLKXOR2X4 U12 ( .A(R[31]), .B(K_sub[46]), .Y(X[46]) );
  CLKXOR2X4 U13 ( .A(R[22]), .B(K_sub[33]), .Y(X[33]) );
  CLKXOR2X4 U14 ( .A(R[16]), .B(K_sub[23]), .Y(X[23]) );
  CLKXOR2X4 U15 ( .A(R[26]), .B(K_sub[39]), .Y(X[39]) );
  CLKXOR2X4 U16 ( .A(R[20]), .B(K_sub[29]), .Y(X[29]) );
  CLKXOR2X2 U17 ( .A(R[4]), .B(K_sub[5]), .Y(X[5]) );
  CLKXOR2X2 U18 ( .A(R[15]), .B(K_sub[22]), .Y(X[22]) );
  CLKXOR2X2 U19 ( .A(R[24]), .B(K_sub[35]), .Y(X[35]) );
  CLKXOR2X2 U20 ( .A(R[21]), .B(K_sub[30]), .Y(X[30]) );
  CLKXOR2X2 U21 ( .A(R[12]), .B(K_sub[17]), .Y(X[17]) );
  CLKXOR2X2 U22 ( .A(R[32]), .B(K_sub[1]), .Y(X[1]) );
  CLKXOR2X2 U23 ( .A(R[13]), .B(K_sub[20]), .Y(X[20]) );
  CLKXOR2X2 U24 ( .A(R[18]), .B(K_sub[27]), .Y(X[27]) );
  CLKXOR2X2 U25 ( .A(R[8]), .B(K_sub[13]), .Y(X[13]) );
  CLKXOR2X2 U26 ( .A(R[4]), .B(K_sub[7]), .Y(X[7]) );
  CLKXOR2X2 U27 ( .A(R[24]), .B(K_sub[37]), .Y(X[37]) );
  CLKXOR2X2 U28 ( .A(R[28]), .B(K_sub[43]), .Y(X[43]) );
  CLKXOR2X2 U29 ( .A(R[1]), .B(K_sub[48]), .Y(X[48]) );
  CLKXOR2X2 U30 ( .A(R[17]), .B(K_sub[24]), .Y(X[24]) );
  CLKXOR2X2 U31 ( .A(R[9]), .B(K_sub[12]), .Y(X[12]) );
  CLKXOR2X2 U32 ( .A(R[13]), .B(K_sub[18]), .Y(X[18]) );
  CLKXOR2X2 U33 ( .A(R[25]), .B(K_sub[36]), .Y(X[36]) );
  XOR2X1 U34 ( .A(R[23]), .B(K_sub[34]), .Y(X[34]) );
  XOR2X1 U35 ( .A(R[9]), .B(K_sub[14]), .Y(X[14]) );
  XOR2X1 U36 ( .A(R[30]), .B(K_sub[45]), .Y(X[45]) );
  XOR2X1 U37 ( .A(R[21]), .B(K_sub[32]), .Y(X[32]) );
  XOR2X1 U38 ( .A(R[25]), .B(K_sub[38]), .Y(X[38]) );
  XOR2X1 U39 ( .A(R[27]), .B(K_sub[40]), .Y(X[40]) );
  XOR2X1 U40 ( .A(R[3]), .B(K_sub[4]), .Y(X[4]) );
  XOR2X1 U41 ( .A(R[11]), .B(K_sub[16]), .Y(X[16]) );
  XOR2X1 U42 ( .A(R[7]), .B(K_sub[10]), .Y(X[10]) );
  XOR2X1 U43 ( .A(R[14]), .B(K_sub[21]), .Y(X[21]) );
  XOR2X1 U44 ( .A(R[6]), .B(K_sub[9]), .Y(X[9]) );
  XOR2X1 U45 ( .A(R[2]), .B(K_sub[3]), .Y(X[3]) );
  XOR2X1 U46 ( .A(R[28]), .B(K_sub[41]), .Y(X[41]) );
  XOR2X1 U47 ( .A(R[17]), .B(K_sub[26]), .Y(X[26]) );
  XOR2X1 U48 ( .A(R[32]), .B(K_sub[47]), .Y(X[47]) );
  XOR2X1 U49 ( .A(R[19]), .B(K_sub[28]), .Y(X[28]) );
endmodule


module sbox1_13 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127;

  OAI222X4 U13 ( .A0(addr[5]), .A1(n101), .B0(n1), .B1(n100), .C0(n99), .C1(n8), .Y(dout[3]) );
  OAI21X2 U42 ( .A0(n4), .A1(n112), .B0(n106), .Y(n123) );
  NAND2X2 U44 ( .A(addr[6]), .B(n13), .Y(n115) );
  NAND2X2 U48 ( .A(addr[1]), .B(n71), .Y(n114) );
  OAI22X2 U49 ( .A0(n72), .A1(n6), .B0(addr[5]), .B1(n120), .Y(n85) );
  NAND2X2 U50 ( .A(n3), .B(n72), .Y(n120) );
  NOR2X2 U51 ( .A(n72), .B(n3), .Y(n124) );
  NOR3X2 U55 ( .A(n2), .B(addr[6]), .C(n8), .Y(n102) );
  NOR2X2 U56 ( .A(n109), .B(n3), .Y(n93) );
  NAND2X2 U57 ( .A(addr[1]), .B(addr[6]), .Y(n109) );
  NAND2X2 U59 ( .A(n13), .B(n71), .Y(n112) );
  NOR2X1 U1 ( .A(n114), .B(n120), .Y(n104) );
  BUFX4 U2 ( .A(addr[4]), .Y(n2) );
  CLKBUFX3 U3 ( .A(addr[2]), .Y(n1) );
  OAI32X1 U4 ( .A0(n112), .A1(n2), .A2(n4), .B0(n115), .B1(n113), .Y(n80) );
  NOR2BXL U5 ( .AN(n118), .B(n1), .Y(n122) );
  CLKBUFX3 U6 ( .A(addr[2]), .Y(n4) );
  INVX3 U7 ( .A(addr[6]), .Y(n71) );
  OAI221X4 U8 ( .A0(addr[5]), .A1(n127), .B0(n126), .B1(n6), .C0(n125), .Y(
        dout[4]) );
  OAI221X4 U9 ( .A0(n88), .A1(n6), .B0(addr[5]), .B1(n87), .C0(n86), .Y(
        dout[2]) );
  OA21XL U10 ( .A0(n95), .A1(n115), .B0(n107), .Y(n119) );
  AOI222XL U11 ( .A0(n12), .A1(n1), .B0(n2), .B1(n110), .C0(n69), .C1(n8), .Y(
        n111) );
  AOI2BB2X1 U12 ( .B0(n2), .B1(n69), .A0N(addr[4]), .A1N(n115), .Y(n91) );
  BUFX4 U14 ( .A(addr[3]), .Y(n3) );
  CLKINVX1 U15 ( .A(n112), .Y(n12) );
  CLKINVX1 U16 ( .A(n113), .Y(n7) );
  NAND2BX1 U17 ( .AN(n104), .B(n119), .Y(n84) );
  CLKXOR2X2 U18 ( .A(n9), .B(n8), .Y(n90) );
  NOR2X1 U19 ( .A(n72), .B(n9), .Y(n118) );
  OAI21XL U20 ( .A0(n9), .A1(n114), .B0(n91), .Y(n92) );
  NAND2X1 U21 ( .A(n93), .B(n72), .Y(n107) );
  NAND2X1 U22 ( .A(n8), .B(n9), .Y(n113) );
  OAI211X1 U23 ( .A0(n72), .A1(n114), .B0(n108), .C0(n107), .Y(n89) );
  CLKINVX1 U24 ( .A(n109), .Y(n69) );
  NAND2X1 U25 ( .A(n124), .B(n11), .Y(n108) );
  CLKINVX1 U26 ( .A(n114), .Y(n70) );
  CLKINVX1 U27 ( .A(n115), .Y(n11) );
  CLKINVX1 U28 ( .A(n95), .Y(n5) );
  AO22X1 U29 ( .A0(n90), .A1(n11), .B0(n9), .B1(n123), .Y(n76) );
  OAI31X1 U30 ( .A0(n8), .A1(n3), .A2(n13), .B0(n103), .Y(n105) );
  AOI31XL U31 ( .A0(n13), .A1(n8), .A2(n2), .B0(n102), .Y(n103) );
  AOI211X1 U32 ( .A0(n10), .A1(n4), .B0(n117), .C0(n116), .Y(n126) );
  CLKINVX1 U33 ( .A(n108), .Y(n10) );
  AOI211X1 U34 ( .A0(n115), .A1(n114), .B0(n113), .C0(n2), .Y(n116) );
  OAI22X1 U35 ( .A0(n120), .A1(n112), .B0(n111), .B1(n9), .Y(n117) );
  AOI211X1 U36 ( .A0(n69), .A1(n118), .B0(n81), .C0(n80), .Y(n88) );
  OAI22X1 U37 ( .A0(n91), .A1(n8), .B0(n3), .B1(n106), .Y(n81) );
  CLKINVX3 U38 ( .A(addr[5]), .Y(n6) );
  NAND2X1 U39 ( .A(n3), .B(n6), .Y(n95) );
  NAND2X1 U40 ( .A(n70), .B(n1), .Y(n106) );
  XOR2X1 U41 ( .A(n82), .B(n2), .Y(n83) );
  NAND2X1 U43 ( .A(n1), .B(n3), .Y(n82) );
  OAI22XL U45 ( .A0(n3), .A1(n13), .B0(n9), .B1(n112), .Y(n94) );
  AOI211XL U46 ( .A0(n98), .A1(n9), .B0(n97), .C0(n104), .Y(n99) );
  OAI22XL U47 ( .A0(n96), .A1(n72), .B0(n95), .B1(n109), .Y(n97) );
  OAI22XL U52 ( .A0(n71), .A1(n6), .B0(n2), .B1(addr[1]), .Y(n98) );
  AOI221XL U53 ( .A0(n5), .A1(addr[6]), .B0(addr[5]), .B1(n94), .C0(n93), .Y(
        n96) );
  OAI21XL U54 ( .A0(addr[1]), .A1(n120), .B0(n119), .Y(n121) );
  AOI221XL U58 ( .A0(n12), .A1(n118), .B0(n93), .B1(n6), .C0(n75), .Y(n78) );
  OAI31X1 U60 ( .A0(n6), .A1(n2), .A2(n74), .B0(n73), .Y(n75) );
  OA21XL U61 ( .A0(n3), .A1(n71), .B0(n109), .Y(n74) );
  OAI21XL U62 ( .A0(n124), .A1(n85), .B0(n70), .Y(n73) );
  OAI21XL U63 ( .A0(n1), .A1(n13), .B0(n109), .Y(n110) );
  INVX4 U64 ( .A(n4), .Y(n8) );
  AOI222XL U65 ( .A0(n124), .A1(n123), .B0(n122), .B1(addr[6]), .C0(n1), .C1(
        n121), .Y(n125) );
  NOR4BBX1 U66 ( .AN(n107), .BN(n106), .C(n105), .D(n104), .Y(n127) );
  AOI222XL U67 ( .A0(n12), .A1(n90), .B0(n89), .B1(n8), .C0(n123), .C1(n72), 
        .Y(n101) );
  AOI2BB2XL U68 ( .B0(addr[5]), .B1(n92), .A0N(n120), .A1N(addr[1]), .Y(n100)
         );
  AOI32X1 U69 ( .A0(n4), .A1(n85), .A2(n12), .B0(n84), .B1(n8), .Y(n86) );
  AOI222XL U70 ( .A0(n124), .A1(n13), .B0(n83), .B1(addr[1]), .C0(n7), .C1(n71), .Y(n87) );
  OAI221X1 U71 ( .A0(n79), .A1(n6), .B0(n4), .B1(n78), .C0(n77), .Y(dout[1])
         );
  AOI32XL U72 ( .A0(addr[6]), .A1(n85), .A2(n1), .B0(n76), .B1(n6), .Y(n77) );
  AOI221X1 U73 ( .A0(n12), .A1(n90), .B0(n4), .B1(n93), .C0(n102), .Y(n79) );
  CLKINVX3 U74 ( .A(n3), .Y(n9) );
  CLKINVX3 U75 ( .A(addr[1]), .Y(n13) );
  CLKINVX3 U76 ( .A(n2), .Y(n72) );
endmodule


module sbox2_13 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147;

  NAND2X2 U55 ( .A(n2), .B(n16), .Y(n136) );
  NAND2X2 U57 ( .A(addr[2]), .B(n5), .Y(n104) );
  NAND2X2 U60 ( .A(addr[5]), .B(addr[2]), .Y(n132) );
  NOR2X2 U61 ( .A(n10), .B(n8), .Y(n101) );
  NAND2X2 U62 ( .A(n83), .B(n9), .Y(n146) );
  NAND2X2 U63 ( .A(n3), .B(n13), .Y(n124) );
  NAND2X2 U64 ( .A(addr[6]), .B(n83), .Y(n122) );
  NAND2X2 U67 ( .A(n3), .B(n2), .Y(n133) );
  AOI222XL U1 ( .A0(n15), .A1(n7), .B0(n88), .B1(n13), .C0(n140), .C1(n8), .Y(
        n89) );
  CLKINVX1 U2 ( .A(n121), .Y(n10) );
  CLKINVX1 U3 ( .A(addr[5]), .Y(n1) );
  INVX3 U4 ( .A(addr[5]), .Y(n5) );
  OAI211X4 U5 ( .A0(n147), .A1(n146), .B0(n145), .C0(n144), .Y(dout[4]) );
  NAND3XL U6 ( .A(n98), .B(n97), .C(n96), .Y(dout[1]) );
  NAND2X1 U7 ( .A(addr[1]), .B(addr[6]), .Y(n121) );
  CLKINVX2 U8 ( .A(addr[1]), .Y(n83) );
  OAI221X1 U9 ( .A0(addr[1]), .A1(n136), .B0(n133), .B1(n83), .C0(n87), .Y(n95) );
  NOR2X1 U10 ( .A(n104), .B(n2), .Y(n141) );
  NOR2X1 U11 ( .A(n124), .B(n2), .Y(n140) );
  CLKBUFX4 U12 ( .A(addr[4]), .Y(n2) );
  NAND2X4 U13 ( .A(addr[1]), .B(n9), .Y(n114) );
  INVX3 U14 ( .A(addr[6]), .Y(n9) );
  NAND2XL U15 ( .A(n102), .B(n16), .Y(n109) );
  AOI211XL U16 ( .A0(n6), .A1(n95), .B0(n94), .C0(n93), .Y(n96) );
  AOI2BB2X1 U17 ( .B0(n5), .B1(n12), .A0N(n104), .A1N(n136), .Y(n117) );
  NOR3BXL U18 ( .AN(n135), .B(n134), .C(n15), .Y(n147) );
  BUFX4 U19 ( .A(addr[3]), .Y(n3) );
  NAND2X1 U20 ( .A(n15), .B(n10), .Y(n113) );
  CLKINVX1 U21 ( .A(n146), .Y(n8) );
  CLKINVX1 U22 ( .A(n115), .Y(n15) );
  CLKINVX1 U23 ( .A(n122), .Y(n11) );
  OAI31X1 U24 ( .A0(n124), .A1(n9), .A2(n5), .B0(n123), .Y(n128) );
  OAI21XL U25 ( .A0(n5), .A1(n83), .B0(n140), .Y(n123) );
  OAI22X1 U26 ( .A0(n122), .A1(n124), .B0(n101), .B1(n132), .Y(n84) );
  INVX1 U27 ( .A(n114), .Y(n7) );
  OAI22X1 U28 ( .A0(n122), .A1(n16), .B0(n82), .B1(n121), .Y(n129) );
  NAND3X1 U29 ( .A(n82), .B(n5), .C(n83), .Y(n111) );
  NAND2X1 U30 ( .A(n16), .B(n82), .Y(n115) );
  OAI21XL U31 ( .A0(n13), .A1(n133), .B0(n135), .Y(n85) );
  OAI22XL U32 ( .A0(n117), .A1(n146), .B0(n116), .B1(n132), .Y(n118) );
  AOI222XL U33 ( .A0(n7), .A1(n115), .B0(n81), .B1(n9), .C0(n15), .C1(n8), .Y(
        n116) );
  CLKINVX1 U34 ( .A(n104), .Y(n4) );
  OAI2BB2XL U35 ( .B0(n114), .B1(n135), .A0N(n126), .A1N(n81), .Y(n106) );
  OAI21XL U36 ( .A0(n112), .A1(n114), .B0(n111), .Y(n120) );
  OAI21XL U37 ( .A0(n133), .A1(n114), .B0(n113), .Y(n119) );
  CLKINVX1 U38 ( .A(n124), .Y(n12) );
  CLKINVX1 U39 ( .A(n136), .Y(n14) );
  CLKINVX1 U40 ( .A(n133), .Y(n81) );
  CLKINVX1 U41 ( .A(n132), .Y(n6) );
  AOI2BB1X1 U42 ( .A0N(n126), .A1N(n125), .B0(n136), .Y(n127) );
  OAI22XL U43 ( .A0(n104), .A1(n114), .B0(n101), .B1(n132), .Y(n102) );
  AO21XL U44 ( .A0(n13), .A1(n14), .B0(n141), .Y(n86) );
  AO21X1 U45 ( .A0(n16), .A1(n4), .B0(n140), .Y(n142) );
  NAND3X1 U46 ( .A(n13), .B(n82), .C(addr[5]), .Y(n135) );
  OAI22X1 U47 ( .A0(addr[5]), .A1(n121), .B0(n122), .B1(n5), .Y(n126) );
  AOI2BB1X1 U48 ( .A0N(n3), .A1N(n1), .B0(n14), .Y(n112) );
  NOR3X1 U49 ( .A(addr[1]), .B(addr[2]), .C(n5), .Y(n125) );
  AOI2BB1XL U50 ( .A0N(n92), .A1N(n91), .B0(addr[5]), .Y(n93) );
  OAI22XL U51 ( .A0(n117), .A1(n114), .B0(n89), .B1(n1), .Y(n94) );
  OAI31XL U52 ( .A0(n114), .A1(n2), .A2(n16), .B0(n90), .Y(n91) );
  OAI21XL U53 ( .A0(n81), .A1(n12), .B0(n11), .Y(n90) );
  NAND2X1 U54 ( .A(n7), .B(n2), .Y(n137) );
  OAI31XL U56 ( .A0(n101), .A1(n3), .A2(addr[2]), .B0(n113), .Y(n92) );
  OAI211X1 U58 ( .A0(n139), .A1(n5), .B0(n138), .C0(n137), .Y(n143) );
  NAND3X1 U59 ( .A(n82), .B(n5), .C(addr[6]), .Y(n138) );
  AOI2BB2X1 U65 ( .B0(n11), .B1(n16), .A0N(n83), .A1N(n136), .Y(n139) );
  OAI22XL U66 ( .A0(addr[5]), .A1(n133), .B0(n3), .B1(n132), .Y(n134) );
  OAI2BB2XL U68 ( .B0(n112), .B1(n122), .A0N(n1), .A1N(n99), .Y(n100) );
  OAI211X1 U69 ( .A0(n146), .A1(n2), .B0(n137), .C0(n113), .Y(n99) );
  NAND3X1 U70 ( .A(n11), .B(n82), .C(n3), .Y(n87) );
  AOI2BB2XL U71 ( .B0(n3), .B1(n105), .A0N(n137), .A1N(n132), .Y(n108) );
  OAI211XL U72 ( .A0(n104), .A1(n146), .B0(n103), .C0(n111), .Y(n105) );
  NAND3XL U73 ( .A(addr[5]), .B(n82), .C(n10), .Y(n103) );
  OAI22XL U74 ( .A0(n3), .A1(n114), .B0(n9), .B1(n115), .Y(n88) );
  NAND4X1 U75 ( .A(n110), .B(n109), .C(n108), .D(n107), .Y(dout[2]) );
  AOI32XL U76 ( .A0(addr[1]), .A1(addr[2]), .A2(n14), .B0(n100), .B1(n13), .Y(
        n110) );
  AOI221XL U77 ( .A0(n125), .A1(addr[4]), .B0(n141), .B1(n11), .C0(n106), .Y(
        n107) );
  AOI33XL U78 ( .A0(n11), .A1(n4), .A2(n2), .B0(n6), .B1(n146), .B2(n3), .Y(
        n145) );
  AOI222XL U79 ( .A0(n143), .A1(n13), .B0(n10), .B1(n142), .C0(n7), .C1(n141), 
        .Y(n144) );
  AOI32XL U80 ( .A0(n4), .A1(n83), .A2(n15), .B0(n8), .B1(n86), .Y(n97) );
  AOI22X1 U81 ( .A0(n10), .A1(n85), .B0(n2), .B1(n84), .Y(n98) );
  NAND2X1 U82 ( .A(n131), .B(n130), .Y(dout[3]) );
  AOI221XL U83 ( .A0(n120), .A1(n13), .B0(addr[2]), .B1(n119), .C0(n118), .Y(
        n131) );
  AOI211X1 U84 ( .A0(n4), .A1(n129), .B0(n128), .C0(n127), .Y(n130) );
  CLKINVX3 U85 ( .A(addr[2]), .Y(n13) );
  CLKINVX3 U86 ( .A(n3), .Y(n16) );
  CLKINVX3 U87 ( .A(n2), .Y(n82) );
endmodule


module sbox3_13 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134;

  NOR2X2 U35 ( .A(n78), .B(addr[3]), .Y(n109) );
  NOR2X2 U50 ( .A(addr[1]), .B(addr[6]), .Y(n108) );
  NOR2X2 U52 ( .A(n11), .B(n3), .Y(n88) );
  NOR2X2 U56 ( .A(n11), .B(n12), .Y(n95) );
  NOR2X1 U1 ( .A(n78), .B(n11), .Y(n107) );
  OAI221X1 U2 ( .A0(n125), .A1(n78), .B0(n4), .B1(addr[1]), .C0(n76), .Y(n105)
         );
  INVXL U3 ( .A(n2), .Y(n1) );
  NOR2X1 U4 ( .A(n17), .B(n4), .Y(n92) );
  NOR2X1 U5 ( .A(n8), .B(n4), .Y(n122) );
  NOR2X1 U6 ( .A(n76), .B(n4), .Y(n96) );
  CLKBUFX3 U7 ( .A(addr[2]), .Y(n4) );
  INVX1 U8 ( .A(addr[2]), .Y(n2) );
  NOR2X1 U9 ( .A(n4), .B(n3), .Y(n111) );
  BUFX4 U10 ( .A(addr[4]), .Y(n3) );
  OAI33X1 U11 ( .A0(n8), .A1(n126), .A2(n12), .B0(n78), .B1(n95), .B2(n120), 
        .Y(n80) );
  INVX3 U12 ( .A(n4), .Y(n12) );
  OAI221X1 U13 ( .A0(addr[5]), .A1(n91), .B0(n90), .B1(n77), .C0(n89), .Y(
        dout[1]) );
  NOR2X4 U14 ( .A(n18), .B(n79), .Y(n125) );
  NOR2X4 U15 ( .A(addr[3]), .B(n3), .Y(n131) );
  NOR2X4 U16 ( .A(n79), .B(addr[6]), .Y(n126) );
  INVX3 U17 ( .A(addr[1]), .Y(n79) );
  NAND2XL U18 ( .A(n95), .B(n125), .Y(n133) );
  OAI211XL U19 ( .A0(n3), .A1(n13), .B0(n129), .C0(n128), .Y(n130) );
  NAND4XL U20 ( .A(n115), .B(n114), .C(n113), .D(n112), .Y(n116) );
  CLKINVX1 U21 ( .A(n133), .Y(n10) );
  INVX1 U22 ( .A(n125), .Y(n15) );
  CLKINVX1 U23 ( .A(n107), .Y(n6) );
  NAND2X1 U24 ( .A(n17), .B(n19), .Y(n123) );
  CLKINVX1 U25 ( .A(n87), .Y(n19) );
  CLKINVX1 U26 ( .A(n121), .Y(n5) );
  CLKINVX1 U27 ( .A(n120), .Y(n16) );
  CLKINVX1 U28 ( .A(n115), .Y(n9) );
  CLKINVX1 U29 ( .A(n108), .Y(n76) );
  NOR2X1 U30 ( .A(n17), .B(n12), .Y(n104) );
  NOR2X1 U31 ( .A(n15), .B(n12), .Y(n110) );
  INVX1 U32 ( .A(n126), .Y(n20) );
  AOI21X1 U33 ( .A0(n11), .A1(n12), .B0(n95), .Y(n121) );
  OAI21XL U34 ( .A0(n111), .A1(n131), .B0(n125), .Y(n83) );
  CLKINVX1 U36 ( .A(n82), .Y(n17) );
  NOR2X1 U37 ( .A(n20), .B(n78), .Y(n87) );
  NOR2X1 U38 ( .A(n125), .B(n108), .Y(n120) );
  OAI21XL U39 ( .A0(n110), .A1(n92), .B0(n131), .Y(n101) );
  NAND2X1 U40 ( .A(n104), .B(n88), .Y(n115) );
  CLKINVX1 U41 ( .A(n88), .Y(n8) );
  CLKINVX1 U42 ( .A(n92), .Y(n13) );
  CLKINVX1 U43 ( .A(n111), .Y(n14) );
  CLKINVX1 U44 ( .A(n122), .Y(n7) );
  OR2X1 U45 ( .A(n104), .B(n96), .Y(n127) );
  OAI221X1 U46 ( .A0(n20), .A1(n14), .B0(n12), .B1(n19), .C0(n94), .Y(n99) );
  AOI221XL U47 ( .A0(n96), .A1(n3), .B0(n93), .B1(n78), .C0(n10), .Y(n94) );
  OAI21XL U48 ( .A0(n12), .A1(n76), .B0(n13), .Y(n93) );
  XNOR2X1 U49 ( .A(addr[5]), .B(addr[3]), .Y(n103) );
  CLKINVX1 U51 ( .A(addr[5]), .Y(n77) );
  OAI221X1 U53 ( .A0(n76), .A1(n14), .B0(n15), .B1(n8), .C0(n106), .Y(n117) );
  AOI221XL U54 ( .A0(addr[3]), .A1(n105), .B0(n104), .B1(n131), .C0(n10), .Y(
        n106) );
  CLKINVX1 U55 ( .A(addr[6]), .Y(n18) );
  NAND3X1 U57 ( .A(n4), .B(n79), .C(n109), .Y(n114) );
  NOR2X1 U58 ( .A(n18), .B(addr[1]), .Y(n82) );
  AOI32XL U59 ( .A0(n12), .A1(n11), .A2(n125), .B0(n124), .B1(n18), .Y(n129)
         );
  AOI22XL U60 ( .A0(n3), .A1(n127), .B0(n126), .B1(n131), .Y(n128) );
  OAI22XL U61 ( .A0(n3), .A1(n2), .B0(n4), .B1(n6), .Y(n124) );
  AOI222XL U62 ( .A0(n111), .A1(n126), .B0(n110), .B1(n11), .C0(n109), .C1(
        n108), .Y(n112) );
  OAI211XL U63 ( .A0(n107), .A1(n131), .B0(n2), .C0(addr[6]), .Y(n113) );
  OAI21XL U64 ( .A0(n1), .A1(addr[1]), .B0(n20), .Y(n81) );
  AOI221XL U65 ( .A0(n87), .A1(n11), .B0(n88), .B1(n126), .C0(n86), .Y(n90) );
  OAI211X1 U66 ( .A0(n85), .A1(n12), .B0(n84), .C0(n83), .Y(n86) );
  AOI222XL U67 ( .A0(n82), .A1(n11), .B0(n108), .B1(n107), .C0(n131), .C1(n79), 
        .Y(n85) );
  OAI21XL U68 ( .A0(n92), .A1(n10), .B0(addr[4]), .Y(n84) );
  AOI221XL U69 ( .A0(n126), .A1(n5), .B0(addr[3]), .B1(n127), .C0(n97), .Y(n98) );
  OAI22X1 U70 ( .A0(n15), .A1(n7), .B0(n6), .B1(n17), .Y(n97) );
  OAI211X1 U71 ( .A0(n76), .A1(n7), .B0(n119), .C0(n118), .Y(dout[3]) );
  AOI32XL U72 ( .A0(n126), .A1(n4), .A2(n103), .B0(n109), .B1(n110), .Y(n119)
         );
  AOI22XL U73 ( .A0(n117), .A1(n77), .B0(addr[5]), .B1(n116), .Y(n118) );
  AOI221XL U74 ( .A0(n122), .A1(n126), .B0(n96), .B1(n109), .C0(n9), .Y(n89)
         );
  AOI221XL U75 ( .A0(n131), .A1(n81), .B0(n95), .B1(n123), .C0(n80), .Y(n91)
         );
  NAND4X1 U76 ( .A(n102), .B(n114), .C(n101), .D(n100), .Y(dout[2]) );
  NAND3XL U77 ( .A(n3), .B(n125), .C(n103), .Y(n102) );
  AOI2BB2XL U78 ( .B0(addr[5]), .B1(n99), .A0N(addr[5]), .A1N(n98), .Y(n100)
         );
  OAI221X1 U79 ( .A0(n134), .A1(n77), .B0(n3), .B1(n133), .C0(n132), .Y(
        dout[4]) );
  AOI32XL U80 ( .A0(n131), .A1(n18), .A2(n1), .B0(n130), .B1(n77), .Y(n132) );
  AOI222XL U81 ( .A0(n5), .A1(n123), .B0(n122), .B1(addr[1]), .C0(n121), .C1(
        n16), .Y(n134) );
  CLKINVX3 U82 ( .A(addr[3]), .Y(n11) );
  CLKINVX3 U83 ( .A(n3), .Y(n78) );
endmodule


module sbox4_13 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126;

  OAI32X4 U12 ( .A0(n6), .A1(n2), .A2(addr[2]), .B0(n5), .B1(n108), .Y(n123)
         );
  OAI222X4 U20 ( .A0(addr[2]), .A1(n92), .B0(n106), .B1(n91), .C0(n90), .C1(
        n72), .Y(dout[2]) );
  OAI222X4 U33 ( .A0(addr[4]), .A1(n106), .B0(n16), .B1(n108), .C0(n2), .C1(
        n118), .Y(n83) );
  NAND2X2 U34 ( .A(addr[4]), .B(n2), .Y(n108) );
  NOR2X2 U43 ( .A(n71), .B(addr[4]), .Y(n113) );
  NOR2X2 U45 ( .A(n5), .B(n2), .Y(n111) );
  NAND2X2 U51 ( .A(n16), .B(n11), .Y(n118) );
  NOR2X2 U52 ( .A(n15), .B(addr[5]), .Y(n97) );
  NAND2X2 U53 ( .A(addr[6]), .B(addr[1]), .Y(n85) );
  NAND2X2 U54 ( .A(addr[1]), .B(n11), .Y(n116) );
  NOR2X2 U55 ( .A(n115), .B(n5), .Y(n121) );
  NAND2X2 U56 ( .A(n71), .B(n15), .Y(n115) );
  NAND2X2 U57 ( .A(addr[5]), .B(n15), .Y(n96) );
  NAND2X2 U58 ( .A(addr[6]), .B(n16), .Y(n106) );
  OAI222X1 U1 ( .A0(n6), .A1(n85), .B0(n97), .B1(n116), .C0(n15), .C1(n118), 
        .Y(n73) );
  CLKINVX1 U2 ( .A(n116), .Y(n10) );
  OAI31X1 U3 ( .A0(n108), .A1(addr[5]), .A2(n12), .B0(n107), .Y(n109) );
  OAI31X4 U4 ( .A0(n118), .A1(n5), .A2(n15), .B0(n117), .Y(n119) );
  CLKINVX1 U5 ( .A(n71), .Y(n1) );
  CLKBUFX3 U6 ( .A(addr[3]), .Y(n2) );
  OAI221X1 U7 ( .A0(addr[2]), .A1(n80), .B0(n118), .B1(n105), .C0(n79), .Y(
        dout[1]) );
  INVX4 U8 ( .A(addr[5]), .Y(n5) );
  AOI222XL U9 ( .A0(n15), .A1(n11), .B0(n113), .B1(n16), .C0(addr[1]), .C1(n71), .Y(n114) );
  OAI222X1 U10 ( .A0(addr[1]), .A1(n84), .B0(n85), .B1(n74), .C0(n71), .C1(
        n107), .Y(n75) );
  NAND2XL U11 ( .A(n1), .B(addr[5]), .Y(n84) );
  AOI211XL U13 ( .A0(n83), .A1(n5), .B0(n82), .C0(n4), .Y(n92) );
  NAND2XL U14 ( .A(n15), .B(n5), .Y(n74) );
  CLKINVX1 U15 ( .A(n118), .Y(n8) );
  CLKINVX1 U16 ( .A(n115), .Y(n14) );
  CLKINVX1 U17 ( .A(n112), .Y(n9) );
  OAI21X1 U18 ( .A0(n10), .A1(n12), .B0(n72), .Y(n112) );
  AOI22X1 U19 ( .A0(n13), .A1(n111), .B0(n12), .B1(n113), .Y(n93) );
  OAI211X1 U21 ( .A0(n16), .A1(n115), .B0(n93), .C0(n3), .Y(n94) );
  CLKINVX1 U22 ( .A(n85), .Y(n13) );
  NAND2X1 U23 ( .A(n97), .B(n71), .Y(n105) );
  NAND2X1 U24 ( .A(n113), .B(n8), .Y(n98) );
  NAND2X1 U25 ( .A(n10), .B(n97), .Y(n107) );
  NAND2X1 U26 ( .A(n118), .B(n85), .Y(n110) );
  OAI21XL U27 ( .A0(n14), .A1(n5), .B0(n108), .Y(n95) );
  CLKINVX1 U28 ( .A(n84), .Y(n7) );
  CLKINVX1 U29 ( .A(addr[2]), .Y(n72) );
  OAI31X1 U30 ( .A0(n15), .A1(addr[6]), .A2(n5), .B0(n87), .Y(n88) );
  OAI21XL U31 ( .A0(n113), .A1(n6), .B0(n13), .Y(n87) );
  OAI211X1 U32 ( .A0(n76), .A1(n15), .B0(n98), .C0(n3), .Y(n77) );
  AOI222XL U35 ( .A0(addr[5]), .A1(addr[6]), .B0(n111), .B1(addr[1]), .C0(n12), 
        .C1(n2), .Y(n76) );
  NAND3XL U36 ( .A(n13), .B(n71), .C(addr[4]), .Y(n117) );
  OAI22XL U37 ( .A0(n116), .A1(n115), .B0(n1), .B1(n112), .Y(n78) );
  CLKINVX3 U38 ( .A(addr[4]), .Y(n15) );
  OAI2BB2XL U39 ( .B0(n115), .B1(n106), .A0N(n5), .A1N(n86), .Y(n89) );
  OAI221XL U40 ( .A0(n116), .A1(addr[4]), .B0(n108), .B1(addr[1]), .C0(n117), 
        .Y(n86) );
  CLKINVX1 U41 ( .A(addr[6]), .Y(n11) );
  CLKINVX1 U42 ( .A(n81), .Y(n4) );
  OAI21XL U44 ( .A0(n96), .A1(n118), .B0(n93), .Y(n82) );
  NAND3X1 U46 ( .A(n101), .B(n100), .C(n99), .Y(n102) );
  AOI32X1 U47 ( .A0(n96), .A1(n71), .A2(n10), .B0(n13), .B1(n95), .Y(n101) );
  AOI2BB2XL U48 ( .B0(n16), .B1(n121), .A0N(n98), .A1N(addr[5]), .Y(n99) );
  OAI21XL U49 ( .A0(n97), .A1(n6), .B0(n12), .Y(n100) );
  AOI2BB2XL U50 ( .B0(n12), .B1(n123), .A0N(n122), .A1N(n72), .Y(n124) );
  AOI211XL U59 ( .A0(n12), .A1(n121), .B0(n120), .C0(n119), .Y(n122) );
  OAI22XL U60 ( .A0(n116), .A1(n115), .B0(addr[5]), .B1(n114), .Y(n120) );
  CLKINVX1 U61 ( .A(n75), .Y(n3) );
  AOI32XL U62 ( .A0(n10), .A1(n96), .A2(n1), .B0(addr[1]), .B1(n121), .Y(n81)
         );
  AOI222XL U63 ( .A0(n12), .A1(n6), .B0(n121), .B1(n116), .C0(n2), .C1(n73), 
        .Y(n80) );
  AOI22XL U64 ( .A0(n78), .A1(n5), .B0(addr[2]), .B1(n77), .Y(n79) );
  NAND2XL U65 ( .A(n111), .B(addr[4]), .Y(n91) );
  AOI211X1 U66 ( .A0(n7), .A1(n110), .B0(n89), .C0(n88), .Y(n90) );
  OAI211X1 U67 ( .A0(n106), .A1(n105), .B0(n104), .C0(n103), .Y(dout[3]) );
  AOI32X1 U68 ( .A0(n2), .A1(n6), .A2(n10), .B0(n94), .B1(n72), .Y(n104) );
  AOI22XL U69 ( .A0(addr[2]), .A1(n102), .B0(n8), .B1(n123), .Y(n103) );
  OAI211X1 U70 ( .A0(addr[2]), .A1(n126), .B0(n125), .C0(n124), .Y(dout[4]) );
  AOI32X1 U71 ( .A0(n13), .A1(n6), .A2(n2), .B0(n9), .B1(n7), .Y(n125) );
  AOI221XL U72 ( .A0(n8), .A1(n111), .B0(n14), .B1(n110), .C0(n109), .Y(n126)
         );
  CLKINVX3 U73 ( .A(n96), .Y(n6) );
  CLKINVX3 U74 ( .A(n106), .Y(n12) );
  CLKINVX3 U75 ( .A(addr[1]), .Y(n16) );
  CLKINVX3 U76 ( .A(n2), .Y(n71) );
endmodule


module sbox5_13 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121;

  OAI222X4 U18 ( .A0(addr[3]), .A1(n106), .B0(n68), .B1(n90), .C0(n70), .C1(n8), .Y(n93) );
  OAI22X2 U40 ( .A0(addr[5]), .A1(n106), .B0(n69), .B1(n114), .Y(n116) );
  NOR2X2 U41 ( .A(n3), .B(addr[3]), .Y(n102) );
  NAND2X2 U45 ( .A(addr[6]), .B(n8), .Y(n114) );
  NAND2X2 U50 ( .A(n8), .B(n68), .Y(n110) );
  NAND2X2 U52 ( .A(addr[1]), .B(n68), .Y(n113) );
  NAND2X2 U54 ( .A(addr[1]), .B(addr[6]), .Y(n106) );
  NAND2X2 U55 ( .A(addr[3]), .B(n70), .Y(n121) );
  CLKINVX1 U1 ( .A(addr[5]), .Y(n1) );
  AOI221XL U2 ( .A0(n93), .A1(n1), .B0(n9), .B1(n13), .C0(n92), .Y(n105) );
  INVX3 U3 ( .A(addr[5]), .Y(n69) );
  OAI221X4 U4 ( .A0(n111), .A1(n110), .B0(n121), .B1(n114), .C0(n109), .Y(n112) );
  OAI221X4 U5 ( .A0(n70), .A1(n114), .B0(n69), .B1(n113), .C0(n120), .Y(n115)
         );
  OAI221X4 U6 ( .A0(n107), .A1(n121), .B0(n111), .B1(n113), .C0(n85), .Y(n86)
         );
  OAI31X1 U7 ( .A0(n14), .A1(addr[5]), .A2(addr[1]), .B0(n81), .Y(n73) );
  OAI32X1 U8 ( .A0(n114), .A1(addr[5]), .A2(n3), .B0(n15), .B1(n107), .Y(n79)
         );
  AOI32XL U9 ( .A0(n13), .A1(n98), .A2(n11), .B0(n2), .B1(n73), .Y(n77) );
  CLKBUFX3 U10 ( .A(addr[4]), .Y(n2) );
  CLKINVX1 U11 ( .A(n81), .Y(n4) );
  NAND2X1 U12 ( .A(n5), .B(n13), .Y(n81) );
  CLKINVX1 U13 ( .A(n110), .Y(n7) );
  CLKXOR2X2 U14 ( .A(n14), .B(n69), .Y(n94) );
  AOI2BB1X1 U15 ( .A0N(n70), .A1N(n1), .B0(n13), .Y(n111) );
  NOR2X1 U16 ( .A(n121), .B(n69), .Y(n91) );
  NOR2BX1 U17 ( .AN(n116), .B(n90), .Y(n83) );
  NAND2X1 U19 ( .A(n7), .B(n69), .Y(n120) );
  CLKINVX1 U20 ( .A(n113), .Y(n11) );
  NAND2X1 U21 ( .A(n11), .B(n69), .Y(n107) );
  CLKINVX1 U22 ( .A(n121), .Y(n15) );
  OAI31X1 U23 ( .A0(n12), .A1(n13), .A2(n113), .B0(n99), .Y(n72) );
  CLKINVX1 U24 ( .A(n106), .Y(n9) );
  OAI2BB2XL U25 ( .B0(n1), .B1(n113), .A0N(n98), .A1N(n5), .Y(n101) );
  CLKINVX1 U26 ( .A(n114), .Y(n5) );
  CLKINVX1 U27 ( .A(n90), .Y(n16) );
  CLKINVX1 U28 ( .A(addr[1]), .Y(n8) );
  CLKINVX1 U29 ( .A(addr[3]), .Y(n14) );
  CLKINVX1 U30 ( .A(addr[6]), .Y(n68) );
  AOI211X1 U31 ( .A0(n91), .A1(addr[1]), .B0(n80), .C0(n79), .Y(n89) );
  OAI2BB2XL U32 ( .B0(n111), .B1(n106), .A0N(n94), .A1N(n7), .Y(n80) );
  AOI211X1 U33 ( .A0(n102), .A1(n84), .B0(n83), .C0(n82), .Y(n85) );
  OAI21XL U34 ( .A0(n68), .A1(n1), .B0(n106), .Y(n84) );
  NOR3XL U35 ( .A(n94), .B(n3), .C(n110), .Y(n82) );
  AOI222XL U36 ( .A0(n9), .A1(n16), .B0(addr[5]), .B1(n108), .C0(n10), .C1(n70), .Y(n109) );
  CLKINVX1 U37 ( .A(n107), .Y(n10) );
  OAI21XL U38 ( .A0(addr[6]), .A1(addr[3]), .B0(n106), .Y(n108) );
  NAND2X1 U39 ( .A(addr[3]), .B(n3), .Y(n90) );
  NAND2X1 U42 ( .A(n2), .B(addr[5]), .Y(n98) );
  NAND2X1 U43 ( .A(n3), .B(n14), .Y(n97) );
  OAI21XL U44 ( .A0(addr[1]), .A1(n97), .B0(n96), .Y(n103) );
  AOI33XL U46 ( .A0(n3), .A1(n95), .A2(addr[5]), .B0(n94), .B1(n70), .B2(
        addr[1]), .Y(n96) );
  OAI21XL U47 ( .A0(n8), .A1(n14), .B0(n114), .Y(n95) );
  OAI21XL U48 ( .A0(addr[6]), .A1(n121), .B0(n99), .Y(n100) );
  NAND2X1 U49 ( .A(n71), .B(n7), .Y(n99) );
  XOR2X1 U51 ( .A(n12), .B(n3), .Y(n71) );
  AOI2BB2XL U53 ( .B0(n102), .B1(n116), .A0N(n2), .A1N(n75), .Y(n76) );
  AOI211X1 U56 ( .A0(n6), .A1(n3), .B0(n74), .C0(n83), .Y(n75) );
  AO22XL U57 ( .A0(n11), .A1(n15), .B0(addr[6]), .B1(n102), .Y(n74) );
  CLKINVX1 U58 ( .A(n120), .Y(n6) );
  CLKINVX1 U59 ( .A(n2), .Y(n12) );
  AO22XL U60 ( .A0(n11), .A1(n16), .B0(addr[6]), .B1(n91), .Y(n92) );
  AOI222XL U61 ( .A0(n116), .A1(n70), .B0(addr[3]), .B1(n115), .C0(n11), .C1(
        n13), .Y(n117) );
  OAI221X1 U62 ( .A0(n2), .A1(n105), .B0(n110), .B1(n121), .C0(n104), .Y(
        dout[3]) );
  AOI222XL U63 ( .A0(n2), .A1(n103), .B0(n102), .B1(n101), .C0(n100), .C1(n1), 
        .Y(n104) );
  OAI211X1 U64 ( .A0(n2), .A1(n89), .B0(n88), .C0(n87), .Y(dout[2]) );
  AOI33XL U65 ( .A0(n15), .A1(n98), .A2(n5), .B0(n3), .B1(n94), .B2(n7), .Y(
        n88) );
  AOI222XL U66 ( .A0(n4), .A1(n69), .B0(n2), .B1(n86), .C0(n91), .C1(n9), .Y(
        n87) );
  OAI211X1 U67 ( .A0(n78), .A1(n69), .B0(n77), .C0(n76), .Y(dout[1]) );
  AOI221XL U68 ( .A0(n15), .A1(addr[1]), .B0(n9), .B1(n13), .C0(n72), .Y(n78)
         );
  OAI211X1 U69 ( .A0(n121), .A1(n120), .B0(n119), .C0(n118), .Y(dout[4]) );
  AOI32XL U70 ( .A0(n13), .A1(n114), .A2(addr[5]), .B0(n2), .B1(n112), .Y(n119) );
  AOI2BB2X1 U71 ( .B0(n4), .B1(n69), .A0N(n2), .A1N(n117), .Y(n118) );
  BUFX4 U72 ( .A(addr[2]), .Y(n3) );
  CLKINVX3 U73 ( .A(n97), .Y(n13) );
  CLKINVX3 U74 ( .A(n3), .Y(n70) );
endmodule


module sbox6_13 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147;

  NAND2X2 U39 ( .A(n138), .B(addr[3]), .Y(n147) );
  NOR2X2 U47 ( .A(n84), .B(n12), .Y(n138) );
  NOR2X2 U50 ( .A(n85), .B(n4), .Y(n119) );
  NOR2X2 U58 ( .A(n81), .B(n85), .Y(n125) );
  NAND2X2 U61 ( .A(n97), .B(n103), .Y(n112) );
  NOR2X2 U62 ( .A(n83), .B(addr[1]), .Y(n103) );
  NOR2X2 U63 ( .A(n81), .B(addr[3]), .Y(n97) );
  NAND2X2 U64 ( .A(n117), .B(n131), .Y(n140) );
  NOR2X2 U65 ( .A(n5), .B(addr[3]), .Y(n131) );
  NOR2X2 U66 ( .A(n13), .B(addr[6]), .Y(n117) );
  NOR2X1 U1 ( .A(n84), .B(addr[3]), .Y(n102) );
  OAI222X1 U2 ( .A0(n91), .A1(n7), .B0(n1), .B1(n18), .C0(addr[5]), .C1(n82), 
        .Y(n92) );
  CLKINVX1 U3 ( .A(n84), .Y(n1) );
  BUFX4 U4 ( .A(addr[2]), .Y(n5) );
  CLKINVX1 U5 ( .A(addr[3]), .Y(n2) );
  OAI22X1 U6 ( .A0(n85), .A1(n83), .B0(addr[1]), .B1(n82), .Y(n142) );
  AOI211X1 U7 ( .A0(n7), .A1(n85), .B0(n131), .C0(n143), .Y(n121) );
  INVX3 U8 ( .A(addr[3]), .Y(n85) );
  CLKINVX1 U9 ( .A(n81), .Y(n3) );
  INVX4 U10 ( .A(n4), .Y(n81) );
  CLKBUFX3 U11 ( .A(addr[4]), .Y(n4) );
  OAI221X1 U12 ( .A0(n83), .A1(n17), .B0(n85), .B1(n10), .C0(n86), .Y(n90) );
  INVX3 U13 ( .A(n96), .Y(n10) );
  OAI221X4 U14 ( .A0(n123), .A1(n15), .B0(n12), .B1(n7), .C0(n9), .Y(n124) );
  NOR2X4 U15 ( .A(addr[1]), .B(addr[6]), .Y(n130) );
  NOR2X4 U16 ( .A(n5), .B(addr[5]), .Y(n143) );
  INVX1 U17 ( .A(n130), .Y(n16) );
  CLKINVX1 U18 ( .A(n125), .Y(n17) );
  NAND2X1 U19 ( .A(n16), .B(n10), .Y(n105) );
  INVXL U20 ( .A(n121), .Y(n6) );
  CLKINVX1 U21 ( .A(n138), .Y(n11) );
  CLKINVX1 U22 ( .A(n117), .Y(n12) );
  CLKINVX1 U23 ( .A(n119), .Y(n82) );
  NOR2X1 U24 ( .A(n10), .B(n123), .Y(n144) );
  NOR2X1 U25 ( .A(n13), .B(n83), .Y(n96) );
  CLKINVX1 U26 ( .A(n103), .Y(n15) );
  OAI211X1 U27 ( .A0(n16), .A1(n17), .B0(n104), .C0(n112), .Y(n108) );
  OAI21XL U28 ( .A0(n103), .A1(n117), .B0(n102), .Y(n104) );
  OAI21XL U29 ( .A0(n132), .A1(n83), .B0(n2), .Y(n86) );
  AOI21X1 U30 ( .A0(n81), .A1(n102), .B0(n125), .Y(n91) );
  OAI2BB2XL U31 ( .B0(n143), .B1(n16), .A0N(n143), .A1N(n117), .Y(n118) );
  CLKINVX1 U32 ( .A(n122), .Y(n9) );
  CLKINVX1 U33 ( .A(n126), .Y(n14) );
  CLKINVX1 U34 ( .A(n97), .Y(n18) );
  NAND2BX1 U35 ( .AN(n144), .B(n137), .Y(n107) );
  CLKINVX1 U36 ( .A(addr[1]), .Y(n13) );
  NOR2X1 U37 ( .A(n10), .B(n1), .Y(n122) );
  NOR2X1 U38 ( .A(addr[1]), .B(n3), .Y(n132) );
  OAI22X1 U40 ( .A0(n82), .A1(n12), .B0(n5), .B1(n14), .Y(n88) );
  NAND2X1 U41 ( .A(n5), .B(n7), .Y(n123) );
  NAND4X1 U42 ( .A(n147), .B(n140), .C(n100), .D(n99), .Y(n101) );
  AOI222XL U43 ( .A0(n98), .A1(n84), .B0(n102), .B1(n130), .C0(n97), .C1(n105), 
        .Y(n99) );
  NAND3X1 U44 ( .A(n5), .B(n82), .C(n96), .Y(n100) );
  OAI221X1 U45 ( .A0(n85), .A1(n15), .B0(n82), .B1(n83), .C0(n14), .Y(n98) );
  AOI22X1 U46 ( .A0(n4), .A1(n115), .B0(addr[5]), .B1(n114), .Y(n129) );
  OAI21XL U48 ( .A0(n121), .A1(n16), .B0(n147), .Y(n115) );
  OAI21XL U49 ( .A0(n113), .A1(n84), .B0(n112), .Y(n114) );
  AOI221XL U51 ( .A0(n119), .A1(n13), .B0(n130), .B1(addr[3]), .C0(n111), .Y(
        n113) );
  OAI22XL U52 ( .A0(n12), .A1(n81), .B0(addr[3]), .B1(n10), .Y(n111) );
  AOI211X1 U53 ( .A0(n4), .A1(n135), .B0(n134), .C0(n133), .Y(n136) );
  OA21XL U54 ( .A0(n2), .A1(n1), .B0(n132), .Y(n133) );
  OAI2BB2XL U55 ( .B0(n3), .B1(n9), .A0N(n131), .A1N(n130), .Y(n134) );
  OAI22X1 U56 ( .A0(n5), .A1(n12), .B0(n84), .B1(n10), .Y(n135) );
  CLKINVX3 U57 ( .A(addr[5]), .Y(n7) );
  AOI2BB2X1 U59 ( .B0(n5), .B1(n130), .A0N(n1), .A1N(n15), .Y(n137) );
  NOR2X1 U60 ( .A(n15), .B(n3), .Y(n126) );
  AOI2BB2XL U67 ( .B0(n143), .B1(n90), .A0N(n89), .A1N(n7), .Y(n94) );
  AOI211X1 U68 ( .A0(n122), .A1(n4), .B0(n88), .C0(n87), .Y(n89) );
  OAI32X1 U69 ( .A0(n15), .A1(n85), .A2(n84), .B0(n11), .B1(n18), .Y(n87) );
  NAND3X1 U70 ( .A(n147), .B(n140), .C(n139), .Y(n141) );
  AOI32X1 U71 ( .A0(n5), .A1(n13), .A2(n4), .B0(n138), .B1(n81), .Y(n139) );
  AO22XL U72 ( .A0(n143), .A1(n3), .B0(n116), .B1(n81), .Y(n120) );
  OAI21XL U73 ( .A0(n1), .A1(n7), .B0(n123), .Y(n116) );
  CLKINVX1 U74 ( .A(n106), .Y(n8) );
  AOI32XL U75 ( .A0(n105), .A1(n81), .A2(n2), .B0(addr[1]), .B1(n125), .Y(n106) );
  OAI211X1 U76 ( .A0(n81), .A1(n140), .B0(n110), .C0(n109), .Y(dout[2]) );
  AOI222XL U77 ( .A0(n108), .A1(n7), .B0(n143), .B1(n8), .C0(n119), .C1(n107), 
        .Y(n109) );
  AOI2BB2XL U78 ( .B0(addr[5]), .B1(n101), .A0N(n84), .A1N(n112), .Y(n110) );
  OAI211X1 U79 ( .A0(n3), .A1(n147), .B0(n146), .C0(n145), .Y(dout[4]) );
  AOI222XL U80 ( .A0(n144), .A1(n85), .B0(n143), .B1(n142), .C0(n141), .C1(n7), 
        .Y(n145) );
  OA22X1 U81 ( .A0(n17), .A1(n137), .B0(n136), .B1(n7), .Y(n146) );
  NAND3X1 U82 ( .A(n129), .B(n128), .C(n127), .Y(dout[3]) );
  AOI32XL U83 ( .A0(n120), .A1(n85), .A2(addr[1]), .B0(n119), .B1(n118), .Y(
        n128) );
  AOI222XL U84 ( .A0(n144), .A1(n81), .B0(n126), .B1(n6), .C0(n125), .C1(n124), 
        .Y(n127) );
  NAND3BX1 U85 ( .AN(n95), .B(n94), .C(n93), .Y(dout[1]) );
  OAI222X1 U86 ( .A0(n140), .A1(n4), .B0(n112), .B1(n84), .C0(n10), .C1(n91), 
        .Y(n95) );
  AOI32XL U87 ( .A0(addr[1]), .A1(n7), .A2(n125), .B0(n130), .B1(n92), .Y(n93)
         );
  CLKINVX3 U88 ( .A(addr[6]), .Y(n83) );
  CLKINVX3 U89 ( .A(n5), .Y(n84) );
endmodule


module sbox7_13 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148;

  OAI222X4 U19 ( .A0(n20), .A1(n129), .B0(n4), .B1(n16), .C0(addr[1]), .C1(n8), 
        .Y(n122) );
  OAI33X4 U33 ( .A0(addr[1]), .A1(n4), .A2(n5), .B0(n17), .B1(n6), .B2(n14), 
        .Y(n97) );
  NOR2X2 U44 ( .A(n84), .B(n4), .Y(n116) );
  NOR2X2 U48 ( .A(addr[1]), .B(addr[6]), .Y(n136) );
  NOR2X2 U51 ( .A(n87), .B(n84), .Y(n125) );
  NOR2X2 U52 ( .A(n17), .B(addr[3]), .Y(n131) );
  NOR2X2 U58 ( .A(n93), .B(n124), .Y(n142) );
  NOR2X2 U60 ( .A(n86), .B(addr[1]), .Y(n93) );
  NOR2X2 U62 ( .A(n12), .B(n3), .Y(n137) );
  NOR2X2 U65 ( .A(n86), .B(n18), .Y(n140) );
  NAND2X1 U1 ( .A(n3), .B(n4), .Y(n119) );
  CLKBUFX3 U2 ( .A(addr[4]), .Y(n4) );
  CLKINVX1 U3 ( .A(n12), .Y(n1) );
  CLKINVX1 U4 ( .A(n6), .Y(n2) );
  CLKBUFX3 U5 ( .A(addr[2]), .Y(n5) );
  OAI22X1 U6 ( .A0(addr[1]), .A1(n8), .B0(n5), .B1(n113), .Y(n100) );
  OAI31X1 U7 ( .A0(n84), .A1(n12), .A2(n18), .B0(n117), .Y(n121) );
  OAI22X1 U8 ( .A0(n4), .A1(n87), .B0(addr[3]), .B1(n11), .Y(n103) );
  NOR2X4 U9 ( .A(n18), .B(addr[6]), .Y(n124) );
  AOI211XL U10 ( .A0(n5), .A1(n15), .B0(n131), .C0(n130), .Y(n132) );
  NOR3XL U11 ( .A(n20), .B(addr[3]), .C(n2), .Y(n130) );
  OAI21XL U12 ( .A0(n3), .A1(n1), .B0(n119), .Y(n89) );
  BUFX4 U13 ( .A(addr[5]), .Y(n3) );
  AOI221XL U14 ( .A0(n140), .A1(n89), .B0(n109), .B1(n15), .C0(n88), .Y(n96)
         );
  CLKINVX1 U15 ( .A(n140), .Y(n17) );
  OAI2BB2XL U16 ( .B0(n142), .B1(n11), .A0N(n141), .A1N(n140), .Y(n143) );
  CLKINVX1 U17 ( .A(n125), .Y(n83) );
  CLKINVX1 U18 ( .A(n142), .Y(n15) );
  NAND2X1 U20 ( .A(n83), .B(n85), .Y(n105) );
  CLKINVX1 U21 ( .A(n123), .Y(n7) );
  CLKINVX1 U22 ( .A(n109), .Y(n10) );
  NAND2X1 U23 ( .A(n124), .B(n84), .Y(n113) );
  CLKINVX1 U24 ( .A(n137), .Y(n11) );
  NOR2X1 U25 ( .A(n11), .B(n84), .Y(n109) );
  CLKINVX1 U26 ( .A(n136), .Y(n20) );
  OAI22XL U27 ( .A0(n137), .A1(n16), .B0(n18), .B1(n10), .Y(n146) );
  OAI21X1 U28 ( .A0(n12), .A1(n83), .B0(n129), .Y(n141) );
  NAND2X1 U29 ( .A(n116), .B(n87), .Y(n129) );
  CLKINVX1 U30 ( .A(n93), .Y(n19) );
  OAI21XL U31 ( .A0(n119), .A1(n19), .B0(n118), .Y(n120) );
  OAI21XL U32 ( .A0(n125), .A1(n137), .B0(n124), .Y(n118) );
  NOR2X1 U34 ( .A(n87), .B(n8), .Y(n123) );
  CLKINVX1 U35 ( .A(n145), .Y(n8) );
  OAI22XL U36 ( .A0(n137), .A1(n113), .B0(n86), .B1(n7), .Y(n88) );
  CLKINVX1 U37 ( .A(n116), .Y(n14) );
  CLKINVX1 U38 ( .A(n131), .Y(n16) );
  CLKINVX1 U39 ( .A(n134), .Y(n85) );
  NOR2XL U40 ( .A(n125), .B(n12), .Y(n110) );
  CLKINVX1 U41 ( .A(n119), .Y(n13) );
  CLKINVX1 U42 ( .A(n103), .Y(n9) );
  OA21XL U43 ( .A0(n21), .A1(n19), .B0(n117), .Y(n102) );
  CLKINVX1 U45 ( .A(n105), .Y(n21) );
  OAI2BB1XL U46 ( .A0N(n103), .A1N(n124), .B0(n102), .Y(n104) );
  OAI22X1 U47 ( .A0(n87), .A1(n14), .B0(n4), .B1(n85), .Y(n112) );
  NOR4X1 U49 ( .A(n4), .B(addr[3]), .C(n18), .D(n6), .Y(n99) );
  XNOR2X1 U50 ( .A(addr[6]), .B(n5), .Y(n101) );
  AOI211X1 U53 ( .A0(n116), .A1(addr[6]), .B0(n115), .C0(n114), .Y(n128) );
  OAI222X1 U54 ( .A0(n111), .A1(n17), .B0(n110), .B1(n19), .C0(n20), .C1(n10), 
        .Y(n115) );
  OAI2BB2XL U55 ( .B0(n13), .B1(n113), .A0N(n18), .A1N(n112), .Y(n114) );
  OA21XL U56 ( .A0(n84), .A1(n3), .B0(n7), .Y(n111) );
  NAND2X1 U57 ( .A(n5), .B(n136), .Y(n133) );
  CLKINVX1 U59 ( .A(addr[6]), .Y(n86) );
  AOI211X1 U61 ( .A0(n131), .A1(n3), .B0(n92), .C0(n91), .Y(n95) );
  OAI221X1 U63 ( .A0(n18), .A1(n8), .B0(n17), .B1(n11), .C0(n102), .Y(n92) );
  OAI31X1 U64 ( .A0(n84), .A1(n12), .A2(n20), .B0(n90), .Y(n91) );
  AO21XL U66 ( .A0(n119), .A1(n129), .B0(addr[6]), .Y(n90) );
  NOR2X1 U67 ( .A(n12), .B(addr[3]), .Y(n145) );
  AOI21XL U68 ( .A0(addr[3]), .A1(n98), .B0(n97), .Y(n108) );
  OAI2BB1XL U69 ( .A0N(n6), .A1N(n124), .B0(n133), .Y(n98) );
  NAND3X1 U70 ( .A(n136), .B(n84), .C(n3), .Y(n117) );
  NOR2X1 U71 ( .A(addr[3]), .B(n3), .Y(n134) );
  OAI21X1 U72 ( .A0(n5), .A1(n142), .B0(n133), .Y(n138) );
  OAI22XL U73 ( .A0(n142), .A1(n14), .B0(n1), .B1(n132), .Y(n135) );
  AO21X1 U74 ( .A0(n139), .A1(n87), .B0(n138), .Y(n144) );
  OAI21XL U75 ( .A0(n2), .A1(n18), .B0(n19), .Y(n139) );
  OAI221X1 U76 ( .A0(n96), .A1(n6), .B0(n5), .B1(n95), .C0(n94), .Y(dout[1])
         );
  AOI2BB2X1 U77 ( .B0(n93), .B1(n112), .A0N(n133), .A1N(n9), .Y(n94) );
  OAI211X1 U78 ( .A0(n128), .A1(n6), .B0(n127), .C0(n126), .Y(dout[3]) );
  AOI32XL U79 ( .A0(n125), .A1(n1), .A2(n124), .B0(n123), .B1(n136), .Y(n126)
         );
  OAI31X1 U80 ( .A0(n122), .A1(n121), .A2(n120), .B0(n6), .Y(n127) );
  OAI221X1 U81 ( .A0(n3), .A1(n108), .B0(n107), .B1(n87), .C0(n106), .Y(
        dout[2]) );
  AOI32XL U82 ( .A0(n105), .A1(n6), .A2(n140), .B0(n2), .B1(n104), .Y(n106) );
  AOI211X1 U83 ( .A0(n101), .A1(n4), .B0(n100), .C0(n99), .Y(n107) );
  NAND2X1 U84 ( .A(n148), .B(n147), .Y(dout[4]) );
  AOI222XL U85 ( .A0(n136), .A1(n141), .B0(n3), .B1(n135), .C0(n134), .C1(n138), .Y(n148) );
  AOI222XL U86 ( .A0(n5), .A1(n146), .B0(n145), .B1(n144), .C0(n143), .C1(n6), 
        .Y(n147) );
  CLKINVX3 U87 ( .A(n5), .Y(n6) );
  CLKINVX3 U88 ( .A(n4), .Y(n12) );
  CLKINVX3 U89 ( .A(addr[1]), .Y(n18) );
  CLKINVX3 U90 ( .A(addr[3]), .Y(n84) );
  CLKINVX3 U91 ( .A(n3), .Y(n87) );
endmodule


module sbox8_13 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132;

  NAND2X2 U41 ( .A(addr[6]), .B(n9), .Y(n131) );
  NAND2X2 U48 ( .A(addr[4]), .B(n6), .Y(n123) );
  NAND2X2 U49 ( .A(n2), .B(n74), .Y(n87) );
  NAND2X2 U50 ( .A(addr[1]), .B(n16), .Y(n124) );
  NAND2X2 U54 ( .A(addr[2]), .B(n14), .Y(n116) );
  NAND2X2 U60 ( .A(addr[6]), .B(addr[1]), .Y(n105) );
  NAND2X2 U61 ( .A(n9), .B(n16), .Y(n108) );
  OAI32X1 U1 ( .A0(n16), .A1(addr[4]), .A2(n92), .B0(n115), .B1(n108), .Y(n96)
         );
  OAI31X1 U2 ( .A0(n123), .A1(addr[6]), .A2(n116), .B0(n109), .Y(n110) );
  OAI221X1 U3 ( .A0(n105), .A1(n87), .B0(addr[4]), .B1(n108), .C0(n86), .Y(n90) );
  NAND2X4 U4 ( .A(addr[4]), .B(n2), .Y(n115) );
  AOI222X1 U5 ( .A0(n88), .A1(addr[2]), .B0(n74), .B1(n15), .C0(n75), .C1(n92), 
        .Y(n114) );
  OAI222X1 U6 ( .A0(addr[2]), .A1(n126), .B0(n6), .B1(n125), .C0(n124), .C1(
        n123), .Y(n127) );
  AOI32XL U7 ( .A0(n12), .A1(n13), .A2(n2), .B0(n8), .B1(n117), .Y(n130) );
  OA21XL U8 ( .A0(n75), .A1(n14), .B0(n121), .Y(n78) );
  INVXL U9 ( .A(n119), .Y(n3) );
  INVX3 U10 ( .A(n2), .Y(n6) );
  BUFX4 U11 ( .A(addr[3]), .Y(n2) );
  CLKBUFX3 U12 ( .A(addr[5]), .Y(n1) );
  CLKINVX1 U13 ( .A(n108), .Y(n8) );
  CLKINVX1 U14 ( .A(n107), .Y(n4) );
  CLKINVX1 U15 ( .A(n93), .Y(n5) );
  NAND2X1 U16 ( .A(n6), .B(n74), .Y(n93) );
  NAND2X1 U17 ( .A(n75), .B(n14), .Y(n121) );
  OAI21XL U18 ( .A0(n115), .A1(n14), .B0(n107), .Y(n77) );
  OAI21X1 U19 ( .A0(n74), .A1(n14), .B0(n123), .Y(n88) );
  OAI31XL U20 ( .A0(n115), .A1(n9), .A2(n116), .B0(n118), .Y(n94) );
  CLKINVX1 U21 ( .A(n131), .Y(n7) );
  NAND2X1 U22 ( .A(n13), .B(n6), .Y(n107) );
  OAI22XL U23 ( .A0(n116), .A1(n123), .B0(n13), .B1(n115), .Y(n117) );
  OAI22XL U24 ( .A0(n123), .A1(n108), .B0(n131), .B1(n93), .Y(n95) );
  OAI2BB2XL U25 ( .B0(n115), .B1(n131), .A0N(n88), .A1N(n11), .Y(n89) );
  AOI211XL U26 ( .A0(n108), .A1(n105), .B0(n74), .C0(n121), .Y(n85) );
  CLKINVX1 U27 ( .A(n124), .Y(n12) );
  OAI22XL U28 ( .A0(n13), .A1(n123), .B0(n78), .B1(n87), .Y(n81) );
  NAND2BX2 U29 ( .AN(n78), .B(n6), .Y(n120) );
  NAND2XL U30 ( .A(n115), .B(n93), .Y(n104) );
  OAI2BB2XL U31 ( .B0(n106), .B1(n105), .A0N(n104), .A1N(n12), .Y(n111) );
  NOR2BXL U32 ( .AN(n123), .B(n103), .Y(n106) );
  NAND3X1 U33 ( .A(n104), .B(n9), .C(n13), .Y(n84) );
  AO21X1 U34 ( .A0(n13), .A1(n11), .B0(n101), .Y(n102) );
  OAI33X1 U35 ( .A0(n16), .A1(n6), .A2(n100), .B0(n75), .B1(n103), .B2(n124), 
        .Y(n101) );
  OA22XL U36 ( .A0(n107), .A1(n131), .B0(n120), .B1(n124), .Y(n98) );
  CLKINVX1 U37 ( .A(n125), .Y(n10) );
  OAI21XL U38 ( .A0(n12), .A1(n7), .B0(addr[4]), .Y(n86) );
  NAND2X1 U39 ( .A(n1), .B(n75), .Y(n100) );
  OAI221X1 U40 ( .A0(n124), .A1(n121), .B0(addr[1]), .B1(n120), .C0(n3), .Y(
        n128) );
  OAI31XL U42 ( .A0(n75), .A1(n9), .A2(n6), .B0(n118), .Y(n119) );
  NAND2X1 U43 ( .A(n11), .B(addr[2]), .Y(n125) );
  NAND4XL U44 ( .A(n7), .B(n1), .C(n2), .D(addr[2]), .Y(n109) );
  NAND3X1 U45 ( .A(n13), .B(n16), .C(n2), .Y(n118) );
  OAI21XL U46 ( .A0(n1), .A1(n87), .B0(n114), .Y(n76) );
  OAI22XL U47 ( .A0(n108), .A1(n120), .B0(n79), .B1(n100), .Y(n80) );
  AOI221XL U51 ( .A0(n7), .A1(n6), .B0(n11), .B1(n2), .C0(n91), .Y(n79) );
  NOR2X1 U52 ( .A(n1), .B(n2), .Y(n103) );
  NOR2X1 U53 ( .A(n87), .B(addr[6]), .Y(n91) );
  NOR2X1 U55 ( .A(n6), .B(n1), .Y(n92) );
  CLKINVX1 U56 ( .A(n100), .Y(n15) );
  OA21XL U57 ( .A0(n1), .A1(n115), .B0(n120), .Y(n132) );
  AOI221XL U58 ( .A0(n8), .A1(n2), .B0(n11), .B1(addr[4]), .C0(n122), .Y(n126)
         );
  OAI22XL U59 ( .A0(n2), .A1(n9), .B0(addr[4]), .B1(n131), .Y(n122) );
  OAI211X1 U62 ( .A0(addr[2]), .A1(n99), .B0(n98), .C0(n97), .Y(dout[2]) );
  AOI221XL U63 ( .A0(addr[2]), .A1(n96), .B0(n1), .B1(n95), .C0(n94), .Y(n97)
         );
  AOI221XL U64 ( .A0(n91), .A1(n1), .B0(n90), .B1(n14), .C0(n89), .Y(n99) );
  OAI211X1 U65 ( .A0(n132), .A1(n131), .B0(n130), .C0(n129), .Y(dout[4]) );
  AOI222XL U66 ( .A0(n128), .A1(n74), .B0(n1), .B1(n127), .C0(n4), .C1(n11), 
        .Y(n129) );
  OAI211X1 U67 ( .A0(addr[1]), .A1(n114), .B0(n113), .C0(n112), .Y(dout[3]) );
  AOI221XL U68 ( .A0(n111), .A1(n75), .B0(n4), .B1(n8), .C0(n110), .Y(n112) );
  AOI2BB2XL U69 ( .B0(n102), .B1(n74), .A0N(n115), .A1N(n125), .Y(n113) );
  NAND4BX1 U70 ( .AN(n85), .B(n84), .C(n83), .D(n82), .Y(dout[1]) );
  AOI221XL U71 ( .A0(n7), .A1(n81), .B0(n5), .B1(n10), .C0(n80), .Y(n82) );
  AOI22X1 U72 ( .A0(n11), .A1(n77), .B0(n12), .B1(n76), .Y(n83) );
  CLKINVX3 U73 ( .A(addr[1]), .Y(n9) );
  CLKINVX3 U74 ( .A(n105), .Y(n11) );
  CLKINVX3 U75 ( .A(n116), .Y(n13) );
  CLKINVX3 U76 ( .A(n1), .Y(n14) );
  CLKINVX3 U77 ( .A(addr[6]), .Y(n16) );
  CLKINVX3 U78 ( .A(addr[4]), .Y(n74) );
  CLKINVX3 U79 ( .A(addr[2]), .Y(n75) );
endmodule


module crp_13 ( P, R, K_sub );
  output [1:32] P;
  input [1:32] R;
  input [1:48] K_sub;
  wire   n1;
  wire   [1:48] X;

  sbox1_13 u0 ( .addr(X[1:6]), .dout({P[9], P[17], P[23], P[31]}) );
  sbox2_13 u1 ( .addr({X[7], n1, X[9:12]}), .dout({P[13], P[28], P[2], P[18]})
         );
  sbox3_13 u2 ( .addr(X[13:18]), .dout({P[24], P[16], P[30], P[6]}) );
  sbox4_13 u3 ( .addr(X[19:24]), .dout({P[26], P[20], P[10], P[1]}) );
  sbox5_13 u4 ( .addr(X[25:30]), .dout({P[8], P[14], P[25], P[3]}) );
  sbox6_13 u5 ( .addr(X[31:36]), .dout({P[4], P[29], P[11], P[19]}) );
  sbox7_13 u6 ( .addr(X[37:42]), .dout({P[32], P[12], P[22], P[7]}) );
  sbox8_13 u7 ( .addr(X[43:48]), .dout({P[5], P[27], P[15], P[21]}) );
  XOR2X1 U1 ( .A(R[1]), .B(K_sub[2]), .Y(X[2]) );
  CLKXOR2X4 U2 ( .A(R[5]), .B(K_sub[6]), .Y(X[6]) );
  CLKXOR2X4 U3 ( .A(R[16]), .B(K_sub[25]), .Y(X[25]) );
  CLKXOR2X4 U4 ( .A(R[29]), .B(K_sub[42]), .Y(X[42]) );
  CLKXOR2X4 U5 ( .A(R[16]), .B(K_sub[23]), .Y(X[23]) );
  CLKXOR2X4 U6 ( .A(R[8]), .B(K_sub[11]), .Y(X[11]) );
  CLKXOR2X4 U7 ( .A(R[22]), .B(K_sub[33]), .Y(X[33]) );
  CLKXOR2X4 U8 ( .A(R[26]), .B(K_sub[39]), .Y(X[39]) );
  CLKXOR2X4 U9 ( .A(R[10]), .B(K_sub[15]), .Y(X[15]) );
  XNOR2X1 U10 ( .A(R[5]), .B(K_sub[8]), .Y(X[8]) );
  INVX3 U11 ( .A(X[8]), .Y(n1) );
  CLKXOR2X4 U12 ( .A(R[20]), .B(K_sub[31]), .Y(X[31]) );
  CLKXOR2X4 U13 ( .A(R[31]), .B(K_sub[46]), .Y(X[46]) );
  CLKXOR2X4 U14 ( .A(R[29]), .B(K_sub[44]), .Y(X[44]) );
  CLKXOR2X4 U15 ( .A(R[12]), .B(K_sub[19]), .Y(X[19]) );
  CLKXOR2X4 U16 ( .A(R[20]), .B(K_sub[29]), .Y(X[29]) );
  CLKXOR2X2 U17 ( .A(R[4]), .B(K_sub[5]), .Y(X[5]) );
  CLKXOR2X2 U18 ( .A(R[15]), .B(K_sub[22]), .Y(X[22]) );
  CLKXOR2X2 U19 ( .A(R[24]), .B(K_sub[35]), .Y(X[35]) );
  CLKXOR2X2 U20 ( .A(R[21]), .B(K_sub[30]), .Y(X[30]) );
  CLKXOR2X2 U21 ( .A(R[12]), .B(K_sub[17]), .Y(X[17]) );
  CLKXOR2X2 U22 ( .A(R[32]), .B(K_sub[1]), .Y(X[1]) );
  CLKXOR2X2 U23 ( .A(R[13]), .B(K_sub[20]), .Y(X[20]) );
  CLKXOR2X2 U24 ( .A(R[18]), .B(K_sub[27]), .Y(X[27]) );
  CLKXOR2X2 U25 ( .A(R[8]), .B(K_sub[13]), .Y(X[13]) );
  CLKXOR2X2 U26 ( .A(R[4]), .B(K_sub[7]), .Y(X[7]) );
  CLKXOR2X2 U27 ( .A(R[24]), .B(K_sub[37]), .Y(X[37]) );
  CLKXOR2X2 U28 ( .A(R[28]), .B(K_sub[43]), .Y(X[43]) );
  CLKXOR2X2 U29 ( .A(R[1]), .B(K_sub[48]), .Y(X[48]) );
  CLKXOR2X2 U30 ( .A(R[17]), .B(K_sub[24]), .Y(X[24]) );
  CLKXOR2X2 U31 ( .A(R[9]), .B(K_sub[12]), .Y(X[12]) );
  CLKXOR2X2 U32 ( .A(R[13]), .B(K_sub[18]), .Y(X[18]) );
  CLKXOR2X2 U33 ( .A(R[25]), .B(K_sub[36]), .Y(X[36]) );
  XOR2X1 U34 ( .A(R[23]), .B(K_sub[34]), .Y(X[34]) );
  XOR2X1 U35 ( .A(R[9]), .B(K_sub[14]), .Y(X[14]) );
  XOR2X1 U36 ( .A(R[30]), .B(K_sub[45]), .Y(X[45]) );
  XOR2X1 U37 ( .A(R[21]), .B(K_sub[32]), .Y(X[32]) );
  XOR2X1 U38 ( .A(R[25]), .B(K_sub[38]), .Y(X[38]) );
  XOR2X1 U39 ( .A(R[27]), .B(K_sub[40]), .Y(X[40]) );
  XOR2X1 U40 ( .A(R[3]), .B(K_sub[4]), .Y(X[4]) );
  XOR2X1 U41 ( .A(R[11]), .B(K_sub[16]), .Y(X[16]) );
  XOR2X1 U42 ( .A(R[7]), .B(K_sub[10]), .Y(X[10]) );
  XOR2X1 U43 ( .A(R[14]), .B(K_sub[21]), .Y(X[21]) );
  XOR2X1 U44 ( .A(R[6]), .B(K_sub[9]), .Y(X[9]) );
  XOR2X1 U45 ( .A(R[2]), .B(K_sub[3]), .Y(X[3]) );
  XOR2X1 U46 ( .A(R[28]), .B(K_sub[41]), .Y(X[41]) );
  XOR2X1 U47 ( .A(R[17]), .B(K_sub[26]), .Y(X[26]) );
  XOR2X1 U48 ( .A(R[32]), .B(K_sub[47]), .Y(X[47]) );
  XOR2X1 U49 ( .A(R[19]), .B(K_sub[28]), .Y(X[28]) );
endmodule


module sbox1_12 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127;

  OAI222X4 U13 ( .A0(addr[5]), .A1(n101), .B0(n1), .B1(n100), .C0(n99), .C1(
        n72), .Y(dout[3]) );
  OAI21X2 U42 ( .A0(n4), .A1(n112), .B0(n106), .Y(n123) );
  NAND2X2 U44 ( .A(addr[6]), .B(n8), .Y(n115) );
  NAND2X2 U48 ( .A(addr[1]), .B(n13), .Y(n114) );
  OAI22X2 U49 ( .A0(n71), .A1(n12), .B0(addr[5]), .B1(n120), .Y(n85) );
  NAND2X2 U50 ( .A(n3), .B(n71), .Y(n120) );
  NOR2X2 U51 ( .A(n71), .B(n3), .Y(n124) );
  NOR3X2 U55 ( .A(n2), .B(addr[6]), .C(n72), .Y(n102) );
  NOR2X2 U56 ( .A(n109), .B(n3), .Y(n93) );
  NAND2X2 U57 ( .A(addr[1]), .B(addr[6]), .Y(n109) );
  NAND2X2 U59 ( .A(n8), .B(n13), .Y(n112) );
  NOR2X1 U1 ( .A(n114), .B(n120), .Y(n104) );
  BUFX4 U2 ( .A(addr[4]), .Y(n2) );
  CLKBUFX3 U3 ( .A(addr[2]), .Y(n1) );
  OAI32X1 U4 ( .A0(n112), .A1(n2), .A2(n4), .B0(n115), .B1(n113), .Y(n80) );
  NOR2BXL U5 ( .AN(n118), .B(n1), .Y(n122) );
  CLKBUFX3 U6 ( .A(addr[2]), .Y(n4) );
  INVX3 U7 ( .A(addr[6]), .Y(n13) );
  OAI221X4 U8 ( .A0(n88), .A1(n12), .B0(addr[5]), .B1(n87), .C0(n86), .Y(
        dout[2]) );
  OAI221X4 U9 ( .A0(addr[5]), .A1(n127), .B0(n126), .B1(n12), .C0(n125), .Y(
        dout[4]) );
  OA21XL U10 ( .A0(n95), .A1(n115), .B0(n107), .Y(n119) );
  AOI222XL U11 ( .A0(n7), .A1(n1), .B0(n2), .B1(n110), .C0(n9), .C1(n72), .Y(
        n111) );
  AOI2BB2X1 U12 ( .B0(n2), .B1(n9), .A0N(addr[4]), .A1N(n115), .Y(n91) );
  BUFX4 U14 ( .A(addr[3]), .Y(n3) );
  CLKINVX1 U15 ( .A(n112), .Y(n7) );
  CLKINVX1 U16 ( .A(n113), .Y(n69) );
  NAND2BX1 U17 ( .AN(n104), .B(n119), .Y(n84) );
  CLKXOR2X2 U18 ( .A(n70), .B(n72), .Y(n90) );
  NOR2X1 U19 ( .A(n71), .B(n70), .Y(n118) );
  OAI21XL U20 ( .A0(n70), .A1(n114), .B0(n91), .Y(n92) );
  NAND2X1 U21 ( .A(n93), .B(n71), .Y(n107) );
  NAND2X1 U22 ( .A(n72), .B(n70), .Y(n113) );
  OAI211X1 U23 ( .A0(n71), .A1(n114), .B0(n108), .C0(n107), .Y(n89) );
  CLKINVX1 U24 ( .A(n109), .Y(n9) );
  NAND2X1 U25 ( .A(n124), .B(n6), .Y(n108) );
  CLKINVX1 U26 ( .A(n114), .Y(n10) );
  CLKINVX1 U27 ( .A(n115), .Y(n6) );
  CLKINVX1 U28 ( .A(n95), .Y(n11) );
  AO22X1 U29 ( .A0(n90), .A1(n6), .B0(n70), .B1(n123), .Y(n76) );
  OAI31X1 U30 ( .A0(n72), .A1(n3), .A2(n8), .B0(n103), .Y(n105) );
  AOI31XL U31 ( .A0(n8), .A1(n72), .A2(n2), .B0(n102), .Y(n103) );
  AOI211X1 U32 ( .A0(n5), .A1(n4), .B0(n117), .C0(n116), .Y(n126) );
  CLKINVX1 U33 ( .A(n108), .Y(n5) );
  AOI211X1 U34 ( .A0(n115), .A1(n114), .B0(n113), .C0(n2), .Y(n116) );
  OAI22X1 U35 ( .A0(n120), .A1(n112), .B0(n111), .B1(n70), .Y(n117) );
  AOI211X1 U36 ( .A0(n9), .A1(n118), .B0(n81), .C0(n80), .Y(n88) );
  OAI22X1 U37 ( .A0(n91), .A1(n72), .B0(n3), .B1(n106), .Y(n81) );
  CLKINVX3 U38 ( .A(addr[5]), .Y(n12) );
  NAND2X1 U39 ( .A(n3), .B(n12), .Y(n95) );
  NAND2X1 U40 ( .A(n10), .B(n1), .Y(n106) );
  XOR2X1 U41 ( .A(n82), .B(n2), .Y(n83) );
  NAND2X1 U43 ( .A(n1), .B(n3), .Y(n82) );
  OAI22XL U45 ( .A0(n3), .A1(n8), .B0(n70), .B1(n112), .Y(n94) );
  AOI211XL U46 ( .A0(n98), .A1(n70), .B0(n97), .C0(n104), .Y(n99) );
  OAI22XL U47 ( .A0(n96), .A1(n71), .B0(n95), .B1(n109), .Y(n97) );
  OAI22XL U52 ( .A0(n13), .A1(n12), .B0(n2), .B1(addr[1]), .Y(n98) );
  AOI221XL U53 ( .A0(n11), .A1(addr[6]), .B0(addr[5]), .B1(n94), .C0(n93), .Y(
        n96) );
  OAI21XL U54 ( .A0(addr[1]), .A1(n120), .B0(n119), .Y(n121) );
  AOI221XL U58 ( .A0(n7), .A1(n118), .B0(n93), .B1(n12), .C0(n75), .Y(n78) );
  OAI31X1 U60 ( .A0(n12), .A1(n2), .A2(n74), .B0(n73), .Y(n75) );
  OA21XL U61 ( .A0(n3), .A1(n13), .B0(n109), .Y(n74) );
  OAI21XL U62 ( .A0(n124), .A1(n85), .B0(n10), .Y(n73) );
  OAI21XL U63 ( .A0(n1), .A1(n8), .B0(n109), .Y(n110) );
  INVX4 U64 ( .A(n4), .Y(n72) );
  AOI222XL U65 ( .A0(n124), .A1(n123), .B0(n122), .B1(addr[6]), .C0(n1), .C1(
        n121), .Y(n125) );
  NOR4BBX1 U66 ( .AN(n107), .BN(n106), .C(n105), .D(n104), .Y(n127) );
  AOI222XL U67 ( .A0(n7), .A1(n90), .B0(n89), .B1(n72), .C0(n123), .C1(n71), 
        .Y(n101) );
  AOI2BB2XL U68 ( .B0(addr[5]), .B1(n92), .A0N(n120), .A1N(addr[1]), .Y(n100)
         );
  AOI32X1 U69 ( .A0(n4), .A1(n85), .A2(n7), .B0(n84), .B1(n72), .Y(n86) );
  AOI222XL U70 ( .A0(n124), .A1(n8), .B0(n83), .B1(addr[1]), .C0(n69), .C1(n13), .Y(n87) );
  OAI221X1 U71 ( .A0(n79), .A1(n12), .B0(n4), .B1(n78), .C0(n77), .Y(dout[1])
         );
  AOI32XL U72 ( .A0(addr[6]), .A1(n85), .A2(n1), .B0(n76), .B1(n12), .Y(n77)
         );
  AOI221X1 U73 ( .A0(n7), .A1(n90), .B0(n4), .B1(n93), .C0(n102), .Y(n79) );
  CLKINVX3 U74 ( .A(addr[1]), .Y(n8) );
  CLKINVX3 U75 ( .A(n3), .Y(n70) );
  CLKINVX3 U76 ( .A(n2), .Y(n71) );
endmodule


module sbox2_12 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147;

  NAND2X2 U55 ( .A(n2), .B(n10), .Y(n136) );
  NAND2X2 U57 ( .A(addr[2]), .B(n82), .Y(n104) );
  NAND2X2 U60 ( .A(addr[5]), .B(addr[2]), .Y(n132) );
  NOR2X2 U61 ( .A(n15), .B(n12), .Y(n101) );
  NAND2X2 U62 ( .A(n14), .B(n83), .Y(n146) );
  NAND2X2 U63 ( .A(n3), .B(n5), .Y(n124) );
  NAND2X2 U64 ( .A(addr[6]), .B(n14), .Y(n122) );
  NAND2X2 U67 ( .A(n3), .B(n2), .Y(n133) );
  AOI222XL U1 ( .A0(n9), .A1(n16), .B0(n88), .B1(n5), .C0(n140), .C1(n12), .Y(
        n89) );
  CLKINVX1 U2 ( .A(n121), .Y(n15) );
  NOR2X1 U3 ( .A(n104), .B(n2), .Y(n141) );
  NOR2X1 U4 ( .A(n124), .B(n2), .Y(n140) );
  CLKBUFX4 U5 ( .A(addr[4]), .Y(n2) );
  CLKINVX1 U6 ( .A(addr[5]), .Y(n1) );
  INVX3 U7 ( .A(addr[5]), .Y(n82) );
  OAI211X4 U8 ( .A0(n147), .A1(n146), .B0(n145), .C0(n144), .Y(dout[4]) );
  NAND3XL U9 ( .A(n98), .B(n97), .C(n96), .Y(dout[1]) );
  NAND2X1 U10 ( .A(addr[1]), .B(addr[6]), .Y(n121) );
  CLKINVX2 U11 ( .A(addr[1]), .Y(n14) );
  OAI221X1 U12 ( .A0(addr[1]), .A1(n136), .B0(n133), .B1(n14), .C0(n87), .Y(
        n95) );
  NAND2X4 U13 ( .A(addr[1]), .B(n83), .Y(n114) );
  INVX3 U14 ( .A(addr[6]), .Y(n83) );
  NAND2XL U15 ( .A(n102), .B(n10), .Y(n109) );
  AOI211XL U16 ( .A0(n6), .A1(n95), .B0(n94), .C0(n93), .Y(n96) );
  AOI2BB2X1 U17 ( .B0(n82), .B1(n4), .A0N(n104), .A1N(n136), .Y(n117) );
  NOR3BXL U18 ( .AN(n135), .B(n134), .C(n9), .Y(n147) );
  BUFX4 U19 ( .A(addr[3]), .Y(n3) );
  NAND2X1 U20 ( .A(n9), .B(n15), .Y(n113) );
  CLKINVX1 U21 ( .A(n146), .Y(n12) );
  CLKINVX1 U22 ( .A(n115), .Y(n9) );
  CLKINVX1 U23 ( .A(n122), .Y(n13) );
  OAI31X1 U24 ( .A0(n124), .A1(n83), .A2(n82), .B0(n123), .Y(n128) );
  OAI21XL U25 ( .A0(n82), .A1(n14), .B0(n140), .Y(n123) );
  OAI22X1 U26 ( .A0(n122), .A1(n124), .B0(n101), .B1(n132), .Y(n84) );
  INVX1 U27 ( .A(n114), .Y(n16) );
  OAI22X1 U28 ( .A0(n122), .A1(n10), .B0(n81), .B1(n121), .Y(n129) );
  NAND3X1 U29 ( .A(n81), .B(n82), .C(n14), .Y(n111) );
  NAND2X1 U30 ( .A(n10), .B(n81), .Y(n115) );
  OAI21XL U31 ( .A0(n5), .A1(n133), .B0(n135), .Y(n85) );
  OAI22XL U32 ( .A0(n117), .A1(n146), .B0(n116), .B1(n132), .Y(n118) );
  AOI222XL U33 ( .A0(n16), .A1(n115), .B0(n11), .B1(n83), .C0(n9), .C1(n12), 
        .Y(n116) );
  CLKINVX1 U34 ( .A(n104), .Y(n7) );
  OAI2BB2XL U35 ( .B0(n114), .B1(n135), .A0N(n126), .A1N(n11), .Y(n106) );
  OAI21XL U36 ( .A0(n112), .A1(n114), .B0(n111), .Y(n120) );
  OAI21XL U37 ( .A0(n133), .A1(n114), .B0(n113), .Y(n119) );
  CLKINVX1 U38 ( .A(n124), .Y(n4) );
  CLKINVX1 U39 ( .A(n136), .Y(n8) );
  CLKINVX1 U40 ( .A(n133), .Y(n11) );
  CLKINVX1 U41 ( .A(n132), .Y(n6) );
  AOI2BB1X1 U42 ( .A0N(n126), .A1N(n125), .B0(n136), .Y(n127) );
  OAI22XL U43 ( .A0(n104), .A1(n114), .B0(n101), .B1(n132), .Y(n102) );
  AO21XL U44 ( .A0(n5), .A1(n8), .B0(n141), .Y(n86) );
  AO21X1 U45 ( .A0(n10), .A1(n7), .B0(n140), .Y(n142) );
  NAND3X1 U46 ( .A(n5), .B(n81), .C(addr[5]), .Y(n135) );
  OAI22X1 U47 ( .A0(addr[5]), .A1(n121), .B0(n122), .B1(n82), .Y(n126) );
  AOI2BB1X1 U48 ( .A0N(n3), .A1N(n1), .B0(n8), .Y(n112) );
  NOR3X1 U49 ( .A(addr[1]), .B(addr[2]), .C(n82), .Y(n125) );
  AOI2BB1XL U50 ( .A0N(n92), .A1N(n91), .B0(addr[5]), .Y(n93) );
  OAI22XL U51 ( .A0(n117), .A1(n114), .B0(n89), .B1(n1), .Y(n94) );
  OAI31XL U52 ( .A0(n114), .A1(n2), .A2(n10), .B0(n90), .Y(n91) );
  OAI21XL U53 ( .A0(n11), .A1(n4), .B0(n13), .Y(n90) );
  NAND2X1 U54 ( .A(n16), .B(n2), .Y(n137) );
  OAI31XL U56 ( .A0(n101), .A1(n3), .A2(addr[2]), .B0(n113), .Y(n92) );
  OAI211X1 U58 ( .A0(n139), .A1(n82), .B0(n138), .C0(n137), .Y(n143) );
  NAND3X1 U59 ( .A(n81), .B(n82), .C(addr[6]), .Y(n138) );
  AOI2BB2X1 U65 ( .B0(n13), .B1(n10), .A0N(n14), .A1N(n136), .Y(n139) );
  OAI22XL U66 ( .A0(addr[5]), .A1(n133), .B0(n3), .B1(n132), .Y(n134) );
  OAI2BB2XL U68 ( .B0(n112), .B1(n122), .A0N(n1), .A1N(n99), .Y(n100) );
  OAI211X1 U69 ( .A0(n146), .A1(n2), .B0(n137), .C0(n113), .Y(n99) );
  NAND3X1 U70 ( .A(n13), .B(n81), .C(n3), .Y(n87) );
  AOI2BB2XL U71 ( .B0(n3), .B1(n105), .A0N(n137), .A1N(n132), .Y(n108) );
  OAI211XL U72 ( .A0(n104), .A1(n146), .B0(n103), .C0(n111), .Y(n105) );
  NAND3XL U73 ( .A(addr[5]), .B(n81), .C(n15), .Y(n103) );
  OAI22XL U74 ( .A0(n3), .A1(n114), .B0(n83), .B1(n115), .Y(n88) );
  NAND4X1 U75 ( .A(n110), .B(n109), .C(n108), .D(n107), .Y(dout[2]) );
  AOI32XL U76 ( .A0(addr[1]), .A1(addr[2]), .A2(n8), .B0(n100), .B1(n5), .Y(
        n110) );
  AOI221XL U77 ( .A0(n125), .A1(addr[4]), .B0(n141), .B1(n13), .C0(n106), .Y(
        n107) );
  AOI33XL U78 ( .A0(n13), .A1(n7), .A2(n2), .B0(n6), .B1(n146), .B2(n3), .Y(
        n145) );
  AOI222XL U79 ( .A0(n143), .A1(n5), .B0(n15), .B1(n142), .C0(n16), .C1(n141), 
        .Y(n144) );
  AOI32XL U80 ( .A0(n7), .A1(n14), .A2(n9), .B0(n12), .B1(n86), .Y(n97) );
  AOI22X1 U81 ( .A0(n15), .A1(n85), .B0(n2), .B1(n84), .Y(n98) );
  NAND2X1 U82 ( .A(n131), .B(n130), .Y(dout[3]) );
  AOI221XL U83 ( .A0(n120), .A1(n5), .B0(addr[2]), .B1(n119), .C0(n118), .Y(
        n131) );
  AOI211X1 U84 ( .A0(n7), .A1(n129), .B0(n128), .C0(n127), .Y(n130) );
  CLKINVX3 U85 ( .A(addr[2]), .Y(n5) );
  CLKINVX3 U86 ( .A(n3), .Y(n10) );
  CLKINVX3 U87 ( .A(n2), .Y(n81) );
endmodule


module sbox3_12 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133;

  NOR2X2 U35 ( .A(n78), .B(addr[3]), .Y(n108) );
  NOR2X2 U50 ( .A(addr[1]), .B(addr[6]), .Y(n107) );
  NOR2X2 U52 ( .A(n20), .B(n2), .Y(n87) );
  NOR2X2 U56 ( .A(n20), .B(n76), .Y(n94) );
  NOR2X1 U1 ( .A(n78), .B(n20), .Y(n106) );
  OAI221X1 U2 ( .A0(n124), .A1(n78), .B0(n3), .B1(addr[1]), .C0(n13), .Y(n104)
         );
  OAI22XL U3 ( .A0(n2), .A1(n76), .B0(n3), .B1(n17), .Y(n123) );
  BUFX4 U4 ( .A(addr[4]), .Y(n2) );
  CLKBUFX3 U5 ( .A(n76), .Y(n1) );
  OAI33X1 U6 ( .A0(n19), .A1(n125), .A2(n76), .B0(n78), .B1(n94), .B2(n119), 
        .Y(n79) );
  INVX3 U7 ( .A(n3), .Y(n76) );
  NOR2X1 U8 ( .A(n12), .B(n3), .Y(n91) );
  NOR2X1 U9 ( .A(n19), .B(n3), .Y(n121) );
  NOR2X1 U10 ( .A(n13), .B(n3), .Y(n95) );
  NOR2X1 U11 ( .A(n3), .B(n2), .Y(n110) );
  CLKBUFX4 U12 ( .A(addr[2]), .Y(n3) );
  OAI221X1 U13 ( .A0(addr[5]), .A1(n90), .B0(n89), .B1(n15), .C0(n88), .Y(
        dout[1]) );
  NOR2X4 U14 ( .A(n14), .B(n9), .Y(n124) );
  NOR2X4 U15 ( .A(addr[3]), .B(n2), .Y(n130) );
  NOR2X4 U16 ( .A(n9), .B(addr[6]), .Y(n125) );
  INVX3 U17 ( .A(addr[1]), .Y(n9) );
  NAND2XL U18 ( .A(n94), .B(n124), .Y(n132) );
  OAI211XL U19 ( .A0(n2), .A1(n11), .B0(n128), .C0(n127), .Y(n129) );
  NAND4XL U20 ( .A(n114), .B(n113), .C(n112), .D(n111), .Y(n115) );
  CLKINVX1 U21 ( .A(n132), .Y(n6) );
  INVX1 U22 ( .A(n124), .Y(n4) );
  CLKINVX1 U23 ( .A(n106), .Y(n17) );
  NAND2X1 U24 ( .A(n12), .B(n7), .Y(n122) );
  CLKINVX1 U25 ( .A(n86), .Y(n7) );
  CLKINVX1 U26 ( .A(n120), .Y(n16) );
  CLKINVX1 U27 ( .A(n119), .Y(n5) );
  CLKINVX1 U28 ( .A(n114), .Y(n10) );
  CLKINVX1 U29 ( .A(n107), .Y(n13) );
  NOR2X1 U30 ( .A(n12), .B(n76), .Y(n103) );
  NOR2X1 U31 ( .A(n4), .B(n76), .Y(n109) );
  INVX1 U32 ( .A(n125), .Y(n8) );
  AOI21X1 U33 ( .A0(n20), .A1(n76), .B0(n94), .Y(n120) );
  OAI21XL U34 ( .A0(n110), .A1(n130), .B0(n124), .Y(n82) );
  CLKINVX1 U36 ( .A(n81), .Y(n12) );
  NOR2X1 U37 ( .A(n8), .B(n78), .Y(n86) );
  NOR2X1 U38 ( .A(n124), .B(n107), .Y(n119) );
  OAI21XL U39 ( .A0(n109), .A1(n91), .B0(n130), .Y(n100) );
  NAND2X1 U40 ( .A(n103), .B(n87), .Y(n114) );
  CLKINVX1 U41 ( .A(n87), .Y(n19) );
  CLKINVX1 U42 ( .A(n91), .Y(n11) );
  CLKINVX1 U43 ( .A(n110), .Y(n77) );
  CLKINVX1 U44 ( .A(n121), .Y(n18) );
  OR2X1 U45 ( .A(n103), .B(n95), .Y(n126) );
  OAI221X1 U46 ( .A0(n8), .A1(n77), .B0(n76), .B1(n7), .C0(n93), .Y(n98) );
  AOI221XL U47 ( .A0(n95), .A1(n2), .B0(n92), .B1(n78), .C0(n6), .Y(n93) );
  OAI21XL U48 ( .A0(n1), .A1(n13), .B0(n11), .Y(n92) );
  XNOR2X1 U49 ( .A(addr[5]), .B(addr[3]), .Y(n102) );
  CLKINVX1 U51 ( .A(addr[5]), .Y(n15) );
  OAI221X1 U53 ( .A0(n13), .A1(n77), .B0(n4), .B1(n19), .C0(n105), .Y(n116) );
  AOI221XL U54 ( .A0(addr[3]), .A1(n104), .B0(n103), .B1(n130), .C0(n6), .Y(
        n105) );
  CLKINVX1 U55 ( .A(addr[6]), .Y(n14) );
  NAND3X1 U57 ( .A(n3), .B(n9), .C(n108), .Y(n113) );
  NOR2X1 U58 ( .A(n14), .B(addr[1]), .Y(n81) );
  AOI32XL U59 ( .A0(n1), .A1(n20), .A2(n124), .B0(n123), .B1(n14), .Y(n128) );
  AOI22XL U60 ( .A0(n2), .A1(n126), .B0(n125), .B1(n130), .Y(n127) );
  AOI222XL U61 ( .A0(n110), .A1(n125), .B0(n109), .B1(n20), .C0(n108), .C1(
        n107), .Y(n111) );
  OAI211XL U62 ( .A0(n106), .A1(n130), .B0(n1), .C0(addr[6]), .Y(n112) );
  OAI21XL U63 ( .A0(n3), .A1(addr[1]), .B0(n8), .Y(n80) );
  AOI221XL U64 ( .A0(n86), .A1(n20), .B0(n87), .B1(n125), .C0(n85), .Y(n89) );
  OAI211X1 U65 ( .A0(n84), .A1(n76), .B0(n83), .C0(n82), .Y(n85) );
  AOI222XL U66 ( .A0(n81), .A1(n20), .B0(n107), .B1(n106), .C0(n130), .C1(n9), 
        .Y(n84) );
  OAI21XL U67 ( .A0(n91), .A1(n6), .B0(addr[4]), .Y(n83) );
  AOI221XL U68 ( .A0(n125), .A1(n16), .B0(addr[3]), .B1(n126), .C0(n96), .Y(
        n97) );
  OAI22X1 U69 ( .A0(n4), .A1(n18), .B0(n17), .B1(n12), .Y(n96) );
  OAI211X1 U70 ( .A0(n13), .A1(n18), .B0(n118), .C0(n117), .Y(dout[3]) );
  AOI32XL U71 ( .A0(n125), .A1(n3), .A2(n102), .B0(n108), .B1(n109), .Y(n118)
         );
  AOI22XL U72 ( .A0(n116), .A1(n15), .B0(addr[5]), .B1(n115), .Y(n117) );
  AOI221XL U73 ( .A0(n121), .A1(n125), .B0(n95), .B1(n108), .C0(n10), .Y(n88)
         );
  AOI221XL U74 ( .A0(n130), .A1(n80), .B0(n94), .B1(n122), .C0(n79), .Y(n90)
         );
  NAND4X1 U75 ( .A(n101), .B(n113), .C(n100), .D(n99), .Y(dout[2]) );
  NAND3XL U76 ( .A(n2), .B(n124), .C(n102), .Y(n101) );
  AOI2BB2XL U77 ( .B0(addr[5]), .B1(n98), .A0N(addr[5]), .A1N(n97), .Y(n99) );
  OAI221X1 U78 ( .A0(n133), .A1(n15), .B0(n2), .B1(n132), .C0(n131), .Y(
        dout[4]) );
  AOI32XL U79 ( .A0(n130), .A1(n14), .A2(addr[2]), .B0(n129), .B1(n15), .Y(
        n131) );
  AOI222XL U80 ( .A0(n16), .A1(n122), .B0(n121), .B1(addr[1]), .C0(n120), .C1(
        n5), .Y(n133) );
  CLKINVX3 U81 ( .A(addr[3]), .Y(n20) );
  CLKINVX3 U82 ( .A(n2), .Y(n78) );
endmodule


module sbox4_12 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126;

  OAI32X4 U12 ( .A0(n71), .A1(n2), .A2(addr[2]), .B0(n16), .B1(n108), .Y(n123)
         );
  OAI222X4 U20 ( .A0(addr[2]), .A1(n92), .B0(n106), .B1(n91), .C0(n90), .C1(
        n14), .Y(dout[2]) );
  OAI222X4 U33 ( .A0(addr[4]), .A1(n106), .B0(n6), .B1(n108), .C0(n2), .C1(
        n118), .Y(n83) );
  NAND2X2 U34 ( .A(addr[4]), .B(n2), .Y(n108) );
  NOR2X2 U43 ( .A(n12), .B(addr[4]), .Y(n113) );
  NOR2X2 U45 ( .A(n16), .B(n2), .Y(n111) );
  NAND2X2 U51 ( .A(n6), .B(n15), .Y(n118) );
  NOR2X2 U52 ( .A(n72), .B(addr[5]), .Y(n97) );
  NAND2X2 U53 ( .A(addr[6]), .B(addr[1]), .Y(n85) );
  NAND2X2 U54 ( .A(addr[1]), .B(n15), .Y(n116) );
  NOR2X2 U55 ( .A(n115), .B(n16), .Y(n121) );
  NAND2X2 U56 ( .A(n12), .B(n72), .Y(n115) );
  NAND2X2 U57 ( .A(addr[5]), .B(n72), .Y(n96) );
  NAND2X2 U58 ( .A(addr[6]), .B(n6), .Y(n106) );
  OAI222X1 U1 ( .A0(n71), .A1(n85), .B0(n97), .B1(n116), .C0(n72), .C1(n118), 
        .Y(n73) );
  CLKINVX1 U2 ( .A(n116), .Y(n9) );
  OAI31X4 U3 ( .A0(n118), .A1(n16), .A2(n72), .B0(n117), .Y(n119) );
  CLKINVX1 U4 ( .A(n12), .Y(n1) );
  CLKBUFX3 U5 ( .A(addr[3]), .Y(n2) );
  OAI221X1 U6 ( .A0(addr[2]), .A1(n80), .B0(n118), .B1(n105), .C0(n79), .Y(
        dout[1]) );
  INVX4 U7 ( .A(addr[5]), .Y(n16) );
  OAI31X1 U8 ( .A0(n108), .A1(addr[5]), .A2(n5), .B0(n107), .Y(n109) );
  AOI222XL U9 ( .A0(n72), .A1(n15), .B0(n113), .B1(n6), .C0(addr[1]), .C1(n12), 
        .Y(n114) );
  OAI222X1 U10 ( .A0(addr[1]), .A1(n84), .B0(n85), .B1(n74), .C0(n12), .C1(
        n107), .Y(n75) );
  NAND2XL U11 ( .A(n1), .B(addr[5]), .Y(n84) );
  AOI211XL U13 ( .A0(n83), .A1(n16), .B0(n82), .C0(n7), .Y(n92) );
  NAND2XL U14 ( .A(n72), .B(n16), .Y(n74) );
  CLKINVX1 U15 ( .A(n118), .Y(n3) );
  CLKINVX1 U16 ( .A(n115), .Y(n11) );
  CLKINVX1 U17 ( .A(n112), .Y(n4) );
  OAI21X1 U18 ( .A0(n9), .A1(n5), .B0(n14), .Y(n112) );
  AOI22X1 U19 ( .A0(n10), .A1(n111), .B0(n5), .B1(n113), .Y(n93) );
  OAI211X1 U21 ( .A0(n6), .A1(n115), .B0(n93), .C0(n8), .Y(n94) );
  CLKINVX1 U22 ( .A(n85), .Y(n10) );
  NAND2X1 U23 ( .A(n97), .B(n12), .Y(n105) );
  NAND2X1 U24 ( .A(n113), .B(n3), .Y(n98) );
  NAND2X1 U25 ( .A(n9), .B(n97), .Y(n107) );
  NAND2X1 U26 ( .A(n118), .B(n85), .Y(n110) );
  OAI21XL U27 ( .A0(n11), .A1(n16), .B0(n108), .Y(n95) );
  CLKINVX1 U28 ( .A(n84), .Y(n13) );
  CLKINVX1 U29 ( .A(addr[2]), .Y(n14) );
  OAI31X1 U30 ( .A0(n72), .A1(addr[6]), .A2(n16), .B0(n87), .Y(n88) );
  OAI21XL U31 ( .A0(n113), .A1(n71), .B0(n10), .Y(n87) );
  OAI211X1 U32 ( .A0(n76), .A1(n72), .B0(n98), .C0(n8), .Y(n77) );
  AOI222XL U35 ( .A0(addr[5]), .A1(addr[6]), .B0(n111), .B1(addr[1]), .C0(n5), 
        .C1(n2), .Y(n76) );
  NAND3XL U36 ( .A(n10), .B(n12), .C(addr[4]), .Y(n117) );
  OAI22XL U37 ( .A0(n116), .A1(n115), .B0(n1), .B1(n112), .Y(n78) );
  CLKINVX3 U38 ( .A(addr[4]), .Y(n72) );
  OAI2BB2XL U39 ( .B0(n115), .B1(n106), .A0N(n16), .A1N(n86), .Y(n89) );
  OAI221XL U40 ( .A0(n116), .A1(addr[4]), .B0(n108), .B1(addr[1]), .C0(n117), 
        .Y(n86) );
  CLKINVX1 U41 ( .A(addr[6]), .Y(n15) );
  CLKINVX1 U42 ( .A(n81), .Y(n7) );
  OAI21XL U44 ( .A0(n96), .A1(n118), .B0(n93), .Y(n82) );
  NAND3X1 U46 ( .A(n101), .B(n100), .C(n99), .Y(n102) );
  AOI32X1 U47 ( .A0(n96), .A1(n12), .A2(n9), .B0(n10), .B1(n95), .Y(n101) );
  AOI2BB2XL U48 ( .B0(n6), .B1(n121), .A0N(n98), .A1N(addr[5]), .Y(n99) );
  OAI21XL U49 ( .A0(n97), .A1(n71), .B0(n5), .Y(n100) );
  AOI2BB2XL U50 ( .B0(n5), .B1(n123), .A0N(n122), .A1N(n14), .Y(n124) );
  AOI211XL U59 ( .A0(n5), .A1(n121), .B0(n120), .C0(n119), .Y(n122) );
  OAI22XL U60 ( .A0(n116), .A1(n115), .B0(addr[5]), .B1(n114), .Y(n120) );
  CLKINVX1 U61 ( .A(n75), .Y(n8) );
  AOI32XL U62 ( .A0(n9), .A1(n96), .A2(n1), .B0(addr[1]), .B1(n121), .Y(n81)
         );
  AOI222XL U63 ( .A0(n5), .A1(n71), .B0(n121), .B1(n116), .C0(n2), .C1(n73), 
        .Y(n80) );
  AOI22XL U64 ( .A0(n78), .A1(n16), .B0(addr[2]), .B1(n77), .Y(n79) );
  NAND2XL U65 ( .A(n111), .B(addr[4]), .Y(n91) );
  AOI211X1 U66 ( .A0(n13), .A1(n110), .B0(n89), .C0(n88), .Y(n90) );
  OAI211X1 U67 ( .A0(n106), .A1(n105), .B0(n104), .C0(n103), .Y(dout[3]) );
  AOI32X1 U68 ( .A0(n2), .A1(n71), .A2(n9), .B0(n94), .B1(n14), .Y(n104) );
  AOI22XL U69 ( .A0(addr[2]), .A1(n102), .B0(n3), .B1(n123), .Y(n103) );
  OAI211X1 U70 ( .A0(addr[2]), .A1(n126), .B0(n125), .C0(n124), .Y(dout[4]) );
  AOI32X1 U71 ( .A0(n10), .A1(n71), .A2(n2), .B0(n4), .B1(n13), .Y(n125) );
  AOI221XL U72 ( .A0(n3), .A1(n111), .B0(n11), .B1(n110), .C0(n109), .Y(n126)
         );
  CLKINVX3 U73 ( .A(n106), .Y(n5) );
  CLKINVX3 U74 ( .A(addr[1]), .Y(n6) );
  CLKINVX3 U75 ( .A(n2), .Y(n12) );
  CLKINVX3 U76 ( .A(n96), .Y(n71) );
endmodule


module sbox5_12 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121;

  OAI222X4 U18 ( .A0(addr[3]), .A1(n106), .B0(n14), .B1(n90), .C0(n69), .C1(
        n68), .Y(n93) );
  OAI22X2 U40 ( .A0(addr[5]), .A1(n106), .B0(n11), .B1(n114), .Y(n116) );
  NOR2X2 U41 ( .A(n3), .B(addr[3]), .Y(n102) );
  NAND2X2 U45 ( .A(addr[6]), .B(n68), .Y(n114) );
  NAND2X2 U50 ( .A(n68), .B(n14), .Y(n110) );
  NAND2X2 U52 ( .A(addr[1]), .B(n14), .Y(n113) );
  NAND2X2 U54 ( .A(addr[1]), .B(addr[6]), .Y(n106) );
  NAND2X2 U55 ( .A(addr[3]), .B(n69), .Y(n121) );
  CLKINVX1 U1 ( .A(addr[5]), .Y(n1) );
  AOI221XL U2 ( .A0(n93), .A1(n1), .B0(n15), .B1(n5), .C0(n92), .Y(n105) );
  INVX3 U3 ( .A(addr[5]), .Y(n11) );
  OAI221X4 U4 ( .A0(n111), .A1(n110), .B0(n121), .B1(n114), .C0(n109), .Y(n112) );
  OAI221X4 U5 ( .A0(n69), .A1(n114), .B0(n11), .B1(n113), .C0(n120), .Y(n115)
         );
  OAI221X4 U6 ( .A0(n107), .A1(n121), .B0(n111), .B1(n113), .C0(n85), .Y(n86)
         );
  OAI31X1 U7 ( .A0(n6), .A1(addr[5]), .A2(addr[1]), .B0(n81), .Y(n73) );
  OAI32X1 U8 ( .A0(n114), .A1(addr[5]), .A2(n3), .B0(n7), .B1(n107), .Y(n79)
         );
  AOI32XL U9 ( .A0(n5), .A1(n98), .A2(n13), .B0(n2), .B1(n73), .Y(n77) );
  CLKBUFX3 U10 ( .A(addr[4]), .Y(n2) );
  CLKINVX1 U11 ( .A(n81), .Y(n4) );
  NAND2X1 U12 ( .A(n16), .B(n5), .Y(n81) );
  CLKINVX1 U13 ( .A(n110), .Y(n12) );
  CLKXOR2X2 U14 ( .A(n6), .B(n11), .Y(n94) );
  AOI2BB1X1 U15 ( .A0N(n69), .A1N(n1), .B0(n5), .Y(n111) );
  NOR2X1 U16 ( .A(n121), .B(n11), .Y(n91) );
  NOR2BX1 U17 ( .AN(n116), .B(n90), .Y(n83) );
  NAND2X1 U19 ( .A(n12), .B(n11), .Y(n120) );
  CLKINVX1 U20 ( .A(n113), .Y(n13) );
  NAND2X1 U21 ( .A(n13), .B(n11), .Y(n107) );
  CLKINVX1 U22 ( .A(n121), .Y(n7) );
  OAI31X1 U23 ( .A0(n70), .A1(n5), .A2(n113), .B0(n99), .Y(n72) );
  CLKINVX1 U24 ( .A(n106), .Y(n15) );
  OAI2BB2XL U25 ( .B0(n1), .B1(n113), .A0N(n98), .A1N(n16), .Y(n101) );
  CLKINVX1 U26 ( .A(n114), .Y(n16) );
  CLKINVX1 U27 ( .A(n90), .Y(n8) );
  CLKINVX1 U28 ( .A(addr[1]), .Y(n68) );
  CLKINVX1 U29 ( .A(addr[3]), .Y(n6) );
  CLKINVX1 U30 ( .A(addr[6]), .Y(n14) );
  AOI211X1 U31 ( .A0(n91), .A1(addr[1]), .B0(n80), .C0(n79), .Y(n89) );
  OAI2BB2XL U32 ( .B0(n111), .B1(n106), .A0N(n94), .A1N(n12), .Y(n80) );
  AOI211X1 U33 ( .A0(n102), .A1(n84), .B0(n83), .C0(n82), .Y(n85) );
  OAI21XL U34 ( .A0(n14), .A1(n1), .B0(n106), .Y(n84) );
  NOR3XL U35 ( .A(n94), .B(n3), .C(n110), .Y(n82) );
  AOI222XL U36 ( .A0(n15), .A1(n8), .B0(addr[5]), .B1(n108), .C0(n9), .C1(n69), 
        .Y(n109) );
  CLKINVX1 U37 ( .A(n107), .Y(n9) );
  OAI21XL U38 ( .A0(addr[6]), .A1(addr[3]), .B0(n106), .Y(n108) );
  NAND2X1 U39 ( .A(addr[3]), .B(n3), .Y(n90) );
  NAND2X1 U42 ( .A(n2), .B(addr[5]), .Y(n98) );
  NAND2X1 U43 ( .A(n3), .B(n6), .Y(n97) );
  OAI21XL U44 ( .A0(addr[1]), .A1(n97), .B0(n96), .Y(n103) );
  AOI33XL U46 ( .A0(n3), .A1(n95), .A2(addr[5]), .B0(n94), .B1(n69), .B2(
        addr[1]), .Y(n96) );
  OAI21XL U47 ( .A0(n68), .A1(n6), .B0(n114), .Y(n95) );
  OAI21XL U48 ( .A0(addr[6]), .A1(n121), .B0(n99), .Y(n100) );
  NAND2X1 U49 ( .A(n71), .B(n12), .Y(n99) );
  XOR2X1 U51 ( .A(n70), .B(n3), .Y(n71) );
  AOI2BB2XL U53 ( .B0(n102), .B1(n116), .A0N(n2), .A1N(n75), .Y(n76) );
  AOI211X1 U56 ( .A0(n10), .A1(n3), .B0(n74), .C0(n83), .Y(n75) );
  AO22XL U57 ( .A0(n13), .A1(n7), .B0(addr[6]), .B1(n102), .Y(n74) );
  CLKINVX1 U58 ( .A(n120), .Y(n10) );
  CLKINVX1 U59 ( .A(n2), .Y(n70) );
  AO22XL U60 ( .A0(n13), .A1(n8), .B0(addr[6]), .B1(n91), .Y(n92) );
  AOI222XL U61 ( .A0(n116), .A1(n69), .B0(addr[3]), .B1(n115), .C0(n13), .C1(
        n5), .Y(n117) );
  OAI221X1 U62 ( .A0(n2), .A1(n105), .B0(n110), .B1(n121), .C0(n104), .Y(
        dout[3]) );
  AOI222XL U63 ( .A0(n2), .A1(n103), .B0(n102), .B1(n101), .C0(n100), .C1(n1), 
        .Y(n104) );
  OAI211X1 U64 ( .A0(n2), .A1(n89), .B0(n88), .C0(n87), .Y(dout[2]) );
  AOI33XL U65 ( .A0(n7), .A1(n98), .A2(n16), .B0(n3), .B1(n94), .B2(n12), .Y(
        n88) );
  AOI222XL U66 ( .A0(n4), .A1(n11), .B0(n2), .B1(n86), .C0(n91), .C1(n15), .Y(
        n87) );
  OAI211X1 U67 ( .A0(n78), .A1(n11), .B0(n77), .C0(n76), .Y(dout[1]) );
  AOI221XL U68 ( .A0(n7), .A1(addr[1]), .B0(n15), .B1(n5), .C0(n72), .Y(n78)
         );
  OAI211X1 U69 ( .A0(n121), .A1(n120), .B0(n119), .C0(n118), .Y(dout[4]) );
  AOI32XL U70 ( .A0(n5), .A1(n114), .A2(addr[5]), .B0(n2), .B1(n112), .Y(n119)
         );
  AOI2BB2X1 U71 ( .B0(n4), .B1(n11), .A0N(n2), .A1N(n117), .Y(n118) );
  BUFX4 U72 ( .A(addr[2]), .Y(n3) );
  CLKINVX3 U73 ( .A(n97), .Y(n5) );
  CLKINVX3 U74 ( .A(n3), .Y(n69) );
endmodule


module sbox6_12 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147;

  NAND2X2 U39 ( .A(n138), .B(addr[3]), .Y(n147) );
  NOR2X2 U47 ( .A(n85), .B(n13), .Y(n138) );
  NOR2X2 U50 ( .A(n18), .B(n4), .Y(n119) );
  NOR2X2 U58 ( .A(n84), .B(n18), .Y(n125) );
  NAND2X2 U61 ( .A(n97), .B(n103), .Y(n112) );
  NOR2X2 U62 ( .A(n11), .B(addr[1]), .Y(n103) );
  NOR2X2 U63 ( .A(n84), .B(addr[3]), .Y(n97) );
  NAND2X2 U64 ( .A(n117), .B(n131), .Y(n140) );
  NOR2X2 U65 ( .A(n5), .B(addr[3]), .Y(n131) );
  NOR2X2 U66 ( .A(n82), .B(addr[6]), .Y(n117) );
  NOR2X1 U1 ( .A(n85), .B(addr[3]), .Y(n102) );
  AOI211X1 U2 ( .A0(n83), .A1(n18), .B0(n131), .C0(n143), .Y(n121) );
  CLKINVX1 U3 ( .A(n84), .Y(n1) );
  INVX4 U4 ( .A(n4), .Y(n84) );
  CLKBUFX3 U5 ( .A(addr[4]), .Y(n4) );
  CLKINVX1 U6 ( .A(n85), .Y(n2) );
  OAI222X1 U7 ( .A0(n91), .A1(n83), .B0(n5), .B1(n81), .C0(addr[5]), .C1(n16), 
        .Y(n92) );
  BUFX4 U8 ( .A(addr[2]), .Y(n5) );
  OAI221X1 U9 ( .A0(n11), .A1(n17), .B0(n18), .B1(n8), .C0(n86), .Y(n90) );
  INVX2 U10 ( .A(n96), .Y(n8) );
  CLKINVX1 U11 ( .A(addr[3]), .Y(n3) );
  INVX3 U12 ( .A(addr[3]), .Y(n18) );
  OAI221X4 U13 ( .A0(n123), .A1(n10), .B0(n13), .B1(n83), .C0(n7), .Y(n124) );
  NOR2X4 U14 ( .A(addr[1]), .B(addr[6]), .Y(n130) );
  NOR2X4 U15 ( .A(n5), .B(addr[5]), .Y(n143) );
  INVX1 U16 ( .A(n130), .Y(n14) );
  CLKINVX1 U17 ( .A(n125), .Y(n17) );
  NAND2X1 U18 ( .A(n14), .B(n8), .Y(n105) );
  INVXL U19 ( .A(n121), .Y(n15) );
  CLKINVX1 U20 ( .A(n138), .Y(n12) );
  CLKINVX1 U21 ( .A(n117), .Y(n13) );
  CLKINVX1 U22 ( .A(n119), .Y(n16) );
  NOR2X1 U23 ( .A(n8), .B(n123), .Y(n144) );
  NOR2X1 U24 ( .A(n82), .B(n11), .Y(n96) );
  CLKINVX1 U25 ( .A(n103), .Y(n10) );
  OAI211X1 U26 ( .A0(n14), .A1(n17), .B0(n104), .C0(n112), .Y(n108) );
  OAI21XL U27 ( .A0(n103), .A1(n117), .B0(n102), .Y(n104) );
  OAI21XL U28 ( .A0(n132), .A1(n11), .B0(n3), .Y(n86) );
  AOI21X1 U29 ( .A0(n84), .A1(n102), .B0(n125), .Y(n91) );
  OAI2BB2XL U30 ( .B0(n143), .B1(n14), .A0N(n143), .A1N(n117), .Y(n118) );
  CLKINVX1 U31 ( .A(n122), .Y(n7) );
  CLKINVX1 U32 ( .A(n126), .Y(n9) );
  CLKINVX1 U33 ( .A(n97), .Y(n81) );
  NAND2BX1 U34 ( .AN(n144), .B(n137), .Y(n107) );
  CLKINVX1 U35 ( .A(addr[1]), .Y(n82) );
  NOR2X1 U36 ( .A(n8), .B(n2), .Y(n122) );
  NOR2X1 U37 ( .A(addr[1]), .B(n1), .Y(n132) );
  OAI22X1 U38 ( .A0(n16), .A1(n13), .B0(n5), .B1(n9), .Y(n88) );
  NAND2X1 U40 ( .A(n2), .B(n83), .Y(n123) );
  NAND4X1 U41 ( .A(n147), .B(n140), .C(n100), .D(n99), .Y(n101) );
  AOI222XL U42 ( .A0(n98), .A1(n85), .B0(n102), .B1(n130), .C0(n97), .C1(n105), 
        .Y(n99) );
  NAND3X1 U43 ( .A(n5), .B(n16), .C(n96), .Y(n100) );
  OAI221X1 U44 ( .A0(n18), .A1(n10), .B0(n16), .B1(n11), .C0(n9), .Y(n98) );
  AOI22X1 U45 ( .A0(n4), .A1(n115), .B0(addr[5]), .B1(n114), .Y(n129) );
  OAI21XL U46 ( .A0(n121), .A1(n14), .B0(n147), .Y(n115) );
  OAI21XL U48 ( .A0(n113), .A1(n85), .B0(n112), .Y(n114) );
  AOI221XL U49 ( .A0(n119), .A1(n82), .B0(n130), .B1(addr[3]), .C0(n111), .Y(
        n113) );
  OAI22XL U51 ( .A0(n13), .A1(n84), .B0(addr[3]), .B1(n8), .Y(n111) );
  OAI22XL U52 ( .A0(n18), .A1(n11), .B0(addr[1]), .B1(n16), .Y(n142) );
  AOI211X1 U53 ( .A0(n4), .A1(n135), .B0(n134), .C0(n133), .Y(n136) );
  OA21XL U54 ( .A0(n3), .A1(n2), .B0(n132), .Y(n133) );
  OAI2BB2XL U55 ( .B0(n1), .B1(n7), .A0N(n131), .A1N(n130), .Y(n134) );
  OAI22X1 U56 ( .A0(n5), .A1(n13), .B0(n85), .B1(n8), .Y(n135) );
  CLKINVX3 U57 ( .A(addr[5]), .Y(n83) );
  AOI2BB2X1 U59 ( .B0(n5), .B1(n130), .A0N(n2), .A1N(n10), .Y(n137) );
  NOR2X1 U60 ( .A(n10), .B(n1), .Y(n126) );
  AOI2BB2XL U67 ( .B0(n143), .B1(n90), .A0N(n89), .A1N(n83), .Y(n94) );
  AOI211X1 U68 ( .A0(n122), .A1(n4), .B0(n88), .C0(n87), .Y(n89) );
  OAI32X1 U69 ( .A0(n10), .A1(n18), .A2(n85), .B0(n12), .B1(n81), .Y(n87) );
  NAND3X1 U70 ( .A(n147), .B(n140), .C(n139), .Y(n141) );
  AOI32X1 U71 ( .A0(n5), .A1(n82), .A2(n4), .B0(n138), .B1(n84), .Y(n139) );
  AO22XL U72 ( .A0(n143), .A1(n1), .B0(n116), .B1(n84), .Y(n120) );
  OAI21XL U73 ( .A0(n2), .A1(n83), .B0(n123), .Y(n116) );
  CLKINVX1 U74 ( .A(n106), .Y(n6) );
  AOI32XL U75 ( .A0(n105), .A1(n84), .A2(n3), .B0(addr[1]), .B1(n125), .Y(n106) );
  OAI211X1 U76 ( .A0(n84), .A1(n140), .B0(n110), .C0(n109), .Y(dout[2]) );
  AOI222XL U77 ( .A0(n108), .A1(n83), .B0(n143), .B1(n6), .C0(n119), .C1(n107), 
        .Y(n109) );
  AOI2BB2XL U78 ( .B0(addr[5]), .B1(n101), .A0N(n85), .A1N(n112), .Y(n110) );
  OAI211X1 U79 ( .A0(n1), .A1(n147), .B0(n146), .C0(n145), .Y(dout[4]) );
  AOI222XL U80 ( .A0(n144), .A1(n18), .B0(n143), .B1(n142), .C0(n141), .C1(n83), .Y(n145) );
  OA22X1 U81 ( .A0(n17), .A1(n137), .B0(n136), .B1(n83), .Y(n146) );
  NAND3X1 U82 ( .A(n129), .B(n128), .C(n127), .Y(dout[3]) );
  AOI32XL U83 ( .A0(n120), .A1(n18), .A2(addr[1]), .B0(n119), .B1(n118), .Y(
        n128) );
  AOI222XL U84 ( .A0(n144), .A1(n84), .B0(n126), .B1(n15), .C0(n125), .C1(n124), .Y(n127) );
  NAND3BX1 U85 ( .AN(n95), .B(n94), .C(n93), .Y(dout[1]) );
  OAI222X1 U86 ( .A0(n140), .A1(n4), .B0(n112), .B1(n85), .C0(n8), .C1(n91), 
        .Y(n95) );
  AOI32XL U87 ( .A0(addr[1]), .A1(n83), .A2(n125), .B0(n130), .B1(n92), .Y(n93) );
  CLKINVX3 U88 ( .A(addr[6]), .Y(n11) );
  CLKINVX3 U89 ( .A(n5), .Y(n85) );
endmodule


module sbox7_12 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148;

  OAI222X4 U19 ( .A0(n11), .A1(n129), .B0(n4), .B1(n7), .C0(addr[1]), .C1(n13), 
        .Y(n122) );
  OAI33X4 U33 ( .A0(addr[1]), .A1(n4), .A2(n5), .B0(n8), .B1(n85), .B2(n19), 
        .Y(n97) );
  NOR2X2 U44 ( .A(n87), .B(n4), .Y(n116) );
  NOR2X2 U48 ( .A(addr[1]), .B(addr[6]), .Y(n136) );
  NOR2X2 U51 ( .A(n83), .B(n87), .Y(n125) );
  NOR2X2 U52 ( .A(n8), .B(addr[3]), .Y(n131) );
  NOR2X2 U58 ( .A(n93), .B(n124), .Y(n142) );
  NOR2X2 U60 ( .A(n86), .B(addr[1]), .Y(n93) );
  NOR2X2 U62 ( .A(n17), .B(n3), .Y(n137) );
  NOR2X2 U65 ( .A(n86), .B(n9), .Y(n140) );
  NAND2X1 U1 ( .A(n3), .B(n4), .Y(n119) );
  CLKBUFX3 U2 ( .A(addr[4]), .Y(n4) );
  CLKINVX1 U3 ( .A(n17), .Y(n1) );
  CLKINVX1 U4 ( .A(n85), .Y(n2) );
  CLKBUFX3 U5 ( .A(addr[2]), .Y(n5) );
  OAI22X1 U6 ( .A0(addr[1]), .A1(n13), .B0(n5), .B1(n113), .Y(n100) );
  OAI31X1 U7 ( .A0(n87), .A1(n17), .A2(n9), .B0(n117), .Y(n121) );
  OAI22X1 U8 ( .A0(n4), .A1(n83), .B0(addr[3]), .B1(n16), .Y(n103) );
  NOR2X4 U9 ( .A(n9), .B(addr[6]), .Y(n124) );
  AOI211XL U10 ( .A0(n5), .A1(n6), .B0(n131), .C0(n130), .Y(n132) );
  NOR3XL U11 ( .A(n11), .B(addr[3]), .C(n2), .Y(n130) );
  OAI21XL U12 ( .A0(n3), .A1(n1), .B0(n119), .Y(n89) );
  BUFX4 U13 ( .A(addr[5]), .Y(n3) );
  AOI221XL U14 ( .A0(n140), .A1(n89), .B0(n109), .B1(n6), .C0(n88), .Y(n96) );
  CLKINVX1 U15 ( .A(n140), .Y(n8) );
  OAI2BB2XL U16 ( .B0(n142), .B1(n16), .A0N(n141), .A1N(n140), .Y(n143) );
  CLKINVX1 U17 ( .A(n125), .Y(n21) );
  CLKINVX1 U18 ( .A(n142), .Y(n6) );
  NAND2X1 U20 ( .A(n21), .B(n84), .Y(n105) );
  CLKINVX1 U21 ( .A(n123), .Y(n12) );
  CLKINVX1 U22 ( .A(n109), .Y(n15) );
  NAND2X1 U23 ( .A(n124), .B(n87), .Y(n113) );
  CLKINVX1 U24 ( .A(n137), .Y(n16) );
  NOR2X1 U25 ( .A(n16), .B(n87), .Y(n109) );
  CLKINVX1 U26 ( .A(n136), .Y(n11) );
  OAI22XL U27 ( .A0(n137), .A1(n7), .B0(n9), .B1(n15), .Y(n146) );
  OAI21X1 U28 ( .A0(n17), .A1(n21), .B0(n129), .Y(n141) );
  NAND2X1 U29 ( .A(n116), .B(n83), .Y(n129) );
  CLKINVX1 U30 ( .A(n93), .Y(n10) );
  OAI21XL U31 ( .A0(n119), .A1(n10), .B0(n118), .Y(n120) );
  OAI21XL U32 ( .A0(n125), .A1(n137), .B0(n124), .Y(n118) );
  NOR2X1 U34 ( .A(n83), .B(n13), .Y(n123) );
  CLKINVX1 U35 ( .A(n145), .Y(n13) );
  OAI22XL U36 ( .A0(n137), .A1(n113), .B0(n86), .B1(n12), .Y(n88) );
  CLKINVX1 U37 ( .A(n116), .Y(n19) );
  CLKINVX1 U38 ( .A(n131), .Y(n7) );
  CLKINVX1 U39 ( .A(n134), .Y(n84) );
  NOR2XL U40 ( .A(n125), .B(n17), .Y(n110) );
  CLKINVX1 U41 ( .A(n119), .Y(n18) );
  CLKINVX1 U42 ( .A(n103), .Y(n14) );
  OA21XL U43 ( .A0(n20), .A1(n10), .B0(n117), .Y(n102) );
  CLKINVX1 U45 ( .A(n105), .Y(n20) );
  OAI2BB1XL U46 ( .A0N(n103), .A1N(n124), .B0(n102), .Y(n104) );
  OAI22X1 U47 ( .A0(n83), .A1(n19), .B0(n4), .B1(n84), .Y(n112) );
  NOR4X1 U49 ( .A(n4), .B(addr[3]), .C(n9), .D(n85), .Y(n99) );
  XNOR2X1 U50 ( .A(addr[6]), .B(n5), .Y(n101) );
  AOI211X1 U53 ( .A0(n116), .A1(addr[6]), .B0(n115), .C0(n114), .Y(n128) );
  OAI222X1 U54 ( .A0(n111), .A1(n8), .B0(n110), .B1(n10), .C0(n11), .C1(n15), 
        .Y(n115) );
  OAI2BB2XL U55 ( .B0(n18), .B1(n113), .A0N(n9), .A1N(n112), .Y(n114) );
  OA21XL U56 ( .A0(n87), .A1(n3), .B0(n12), .Y(n111) );
  NAND2X1 U57 ( .A(n5), .B(n136), .Y(n133) );
  CLKINVX1 U59 ( .A(addr[6]), .Y(n86) );
  AOI211X1 U61 ( .A0(n131), .A1(n3), .B0(n92), .C0(n91), .Y(n95) );
  OAI221X1 U63 ( .A0(n9), .A1(n13), .B0(n8), .B1(n16), .C0(n102), .Y(n92) );
  OAI31X1 U64 ( .A0(n87), .A1(n17), .A2(n11), .B0(n90), .Y(n91) );
  AO21XL U66 ( .A0(n119), .A1(n129), .B0(addr[6]), .Y(n90) );
  NOR2X1 U67 ( .A(n17), .B(addr[3]), .Y(n145) );
  AOI21XL U68 ( .A0(addr[3]), .A1(n98), .B0(n97), .Y(n108) );
  OAI2BB1XL U69 ( .A0N(n85), .A1N(n124), .B0(n133), .Y(n98) );
  NAND3X1 U70 ( .A(n136), .B(n87), .C(n3), .Y(n117) );
  NOR2X1 U71 ( .A(addr[3]), .B(n3), .Y(n134) );
  OAI21X1 U72 ( .A0(n5), .A1(n142), .B0(n133), .Y(n138) );
  OAI22XL U73 ( .A0(n142), .A1(n19), .B0(n1), .B1(n132), .Y(n135) );
  AO21X1 U74 ( .A0(n139), .A1(n83), .B0(n138), .Y(n144) );
  OAI21XL U75 ( .A0(n2), .A1(n9), .B0(n10), .Y(n139) );
  OAI221X1 U76 ( .A0(n96), .A1(n85), .B0(n5), .B1(n95), .C0(n94), .Y(dout[1])
         );
  AOI2BB2X1 U77 ( .B0(n93), .B1(n112), .A0N(n133), .A1N(n14), .Y(n94) );
  OAI211X1 U78 ( .A0(n128), .A1(n85), .B0(n127), .C0(n126), .Y(dout[3]) );
  AOI32XL U79 ( .A0(n125), .A1(n1), .A2(n124), .B0(n123), .B1(n136), .Y(n126)
         );
  OAI31X1 U80 ( .A0(n122), .A1(n121), .A2(n120), .B0(n85), .Y(n127) );
  OAI221X1 U81 ( .A0(n3), .A1(n108), .B0(n107), .B1(n83), .C0(n106), .Y(
        dout[2]) );
  AOI32XL U82 ( .A0(n105), .A1(n85), .A2(n140), .B0(n2), .B1(n104), .Y(n106)
         );
  AOI211X1 U83 ( .A0(n101), .A1(n4), .B0(n100), .C0(n99), .Y(n107) );
  NAND2X1 U84 ( .A(n148), .B(n147), .Y(dout[4]) );
  AOI222XL U85 ( .A0(n136), .A1(n141), .B0(n3), .B1(n135), .C0(n134), .C1(n138), .Y(n148) );
  AOI222XL U86 ( .A0(n5), .A1(n146), .B0(n145), .B1(n144), .C0(n143), .C1(n85), 
        .Y(n147) );
  CLKINVX3 U87 ( .A(addr[1]), .Y(n9) );
  CLKINVX3 U88 ( .A(n4), .Y(n17) );
  CLKINVX3 U89 ( .A(n3), .Y(n83) );
  CLKINVX3 U90 ( .A(n5), .Y(n85) );
  CLKINVX3 U91 ( .A(addr[3]), .Y(n87) );
endmodule


module sbox8_12 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132;

  NAND2X2 U41 ( .A(addr[6]), .B(n14), .Y(n131) );
  NAND2X2 U48 ( .A(addr[4]), .B(n7), .Y(n123) );
  NAND2X2 U49 ( .A(n2), .B(n4), .Y(n87) );
  NAND2X2 U50 ( .A(addr[1]), .B(n75), .Y(n124) );
  NAND2X2 U54 ( .A(addr[2]), .B(n74), .Y(n116) );
  NAND2X2 U60 ( .A(addr[6]), .B(addr[1]), .Y(n105) );
  NAND2X2 U61 ( .A(n14), .B(n75), .Y(n108) );
  OAI31X1 U1 ( .A0(n123), .A1(addr[6]), .A2(n116), .B0(n109), .Y(n110) );
  AOI222X1 U2 ( .A0(n88), .A1(addr[2]), .B0(n4), .B1(n8), .C0(n9), .C1(n92), 
        .Y(n114) );
  OAI222X1 U3 ( .A0(addr[2]), .A1(n126), .B0(n7), .B1(n125), .C0(n124), .C1(
        n123), .Y(n127) );
  NAND2X4 U4 ( .A(addr[4]), .B(n2), .Y(n115) );
  OAI32X1 U5 ( .A0(n75), .A1(addr[4]), .A2(n92), .B0(n115), .B1(n108), .Y(n96)
         );
  OAI221X1 U6 ( .A0(n105), .A1(n87), .B0(addr[4]), .B1(n108), .C0(n86), .Y(n90) );
  AOI32XL U7 ( .A0(n16), .A1(n10), .A2(n2), .B0(n13), .B1(n117), .Y(n130) );
  OA21XL U8 ( .A0(n9), .A1(n74), .B0(n121), .Y(n78) );
  INVXL U9 ( .A(n119), .Y(n5) );
  INVX3 U10 ( .A(n2), .Y(n7) );
  BUFX4 U11 ( .A(addr[3]), .Y(n2) );
  CLKBUFX3 U12 ( .A(addr[5]), .Y(n1) );
  CLKINVX1 U13 ( .A(n108), .Y(n13) );
  CLKINVX1 U14 ( .A(n107), .Y(n6) );
  CLKINVX1 U15 ( .A(n93), .Y(n3) );
  NAND2X1 U16 ( .A(n7), .B(n4), .Y(n93) );
  NAND2X1 U17 ( .A(n9), .B(n74), .Y(n121) );
  OAI21XL U18 ( .A0(n115), .A1(n74), .B0(n107), .Y(n77) );
  OAI21X1 U19 ( .A0(n4), .A1(n74), .B0(n123), .Y(n88) );
  OAI31XL U20 ( .A0(n115), .A1(n14), .A2(n116), .B0(n118), .Y(n94) );
  CLKINVX1 U21 ( .A(n131), .Y(n12) );
  NAND2X1 U22 ( .A(n10), .B(n7), .Y(n107) );
  OAI22XL U23 ( .A0(n116), .A1(n123), .B0(n10), .B1(n115), .Y(n117) );
  OAI22XL U24 ( .A0(n123), .A1(n108), .B0(n131), .B1(n93), .Y(n95) );
  OAI2BB2XL U25 ( .B0(n115), .B1(n131), .A0N(n88), .A1N(n15), .Y(n89) );
  AOI211XL U26 ( .A0(n108), .A1(n105), .B0(n4), .C0(n121), .Y(n85) );
  CLKINVX1 U27 ( .A(n124), .Y(n16) );
  OAI22XL U28 ( .A0(n10), .A1(n123), .B0(n78), .B1(n87), .Y(n81) );
  NAND2BX2 U29 ( .AN(n78), .B(n7), .Y(n120) );
  NAND2XL U30 ( .A(n115), .B(n93), .Y(n104) );
  OAI2BB2XL U31 ( .B0(n106), .B1(n105), .A0N(n104), .A1N(n16), .Y(n111) );
  NOR2BXL U32 ( .AN(n123), .B(n103), .Y(n106) );
  NAND3X1 U33 ( .A(n104), .B(n14), .C(n10), .Y(n84) );
  AO21X1 U34 ( .A0(n10), .A1(n15), .B0(n101), .Y(n102) );
  OAI33X1 U35 ( .A0(n75), .A1(n7), .A2(n100), .B0(n9), .B1(n103), .B2(n124), 
        .Y(n101) );
  OA22XL U36 ( .A0(n107), .A1(n131), .B0(n120), .B1(n124), .Y(n98) );
  CLKINVX1 U37 ( .A(n125), .Y(n11) );
  OAI21XL U38 ( .A0(n16), .A1(n12), .B0(addr[4]), .Y(n86) );
  NAND2X1 U39 ( .A(n1), .B(n9), .Y(n100) );
  OAI221X1 U40 ( .A0(n124), .A1(n121), .B0(addr[1]), .B1(n120), .C0(n5), .Y(
        n128) );
  OAI31XL U42 ( .A0(n9), .A1(n14), .A2(n7), .B0(n118), .Y(n119) );
  NAND2X1 U43 ( .A(n15), .B(addr[2]), .Y(n125) );
  NAND4XL U44 ( .A(n12), .B(n1), .C(n2), .D(addr[2]), .Y(n109) );
  NAND3X1 U45 ( .A(n10), .B(n75), .C(n2), .Y(n118) );
  OAI21XL U46 ( .A0(n1), .A1(n87), .B0(n114), .Y(n76) );
  OAI22XL U47 ( .A0(n108), .A1(n120), .B0(n79), .B1(n100), .Y(n80) );
  AOI221XL U51 ( .A0(n12), .A1(n7), .B0(n15), .B1(n2), .C0(n91), .Y(n79) );
  NOR2X1 U52 ( .A(n1), .B(n2), .Y(n103) );
  NOR2X1 U53 ( .A(n87), .B(addr[6]), .Y(n91) );
  NOR2X1 U55 ( .A(n7), .B(n1), .Y(n92) );
  CLKINVX1 U56 ( .A(n100), .Y(n8) );
  OA21XL U57 ( .A0(n1), .A1(n115), .B0(n120), .Y(n132) );
  AOI221XL U58 ( .A0(n13), .A1(n2), .B0(n15), .B1(addr[4]), .C0(n122), .Y(n126) );
  OAI22XL U59 ( .A0(n2), .A1(n14), .B0(addr[4]), .B1(n131), .Y(n122) );
  OAI211X1 U62 ( .A0(addr[2]), .A1(n99), .B0(n98), .C0(n97), .Y(dout[2]) );
  AOI221XL U63 ( .A0(addr[2]), .A1(n96), .B0(n1), .B1(n95), .C0(n94), .Y(n97)
         );
  AOI221XL U64 ( .A0(n91), .A1(n1), .B0(n90), .B1(n74), .C0(n89), .Y(n99) );
  OAI211X1 U65 ( .A0(n132), .A1(n131), .B0(n130), .C0(n129), .Y(dout[4]) );
  AOI222XL U66 ( .A0(n128), .A1(n4), .B0(n1), .B1(n127), .C0(n6), .C1(n15), 
        .Y(n129) );
  OAI211X1 U67 ( .A0(addr[1]), .A1(n114), .B0(n113), .C0(n112), .Y(dout[3]) );
  AOI221XL U68 ( .A0(n111), .A1(n9), .B0(n6), .B1(n13), .C0(n110), .Y(n112) );
  AOI2BB2XL U69 ( .B0(n102), .B1(n4), .A0N(n115), .A1N(n125), .Y(n113) );
  NAND4BX1 U70 ( .AN(n85), .B(n84), .C(n83), .D(n82), .Y(dout[1]) );
  AOI221XL U71 ( .A0(n12), .A1(n81), .B0(n3), .B1(n11), .C0(n80), .Y(n82) );
  AOI22X1 U72 ( .A0(n15), .A1(n77), .B0(n16), .B1(n76), .Y(n83) );
  CLKINVX3 U73 ( .A(addr[4]), .Y(n4) );
  CLKINVX3 U74 ( .A(addr[2]), .Y(n9) );
  CLKINVX3 U75 ( .A(n116), .Y(n10) );
  CLKINVX3 U76 ( .A(addr[1]), .Y(n14) );
  CLKINVX3 U77 ( .A(n105), .Y(n15) );
  CLKINVX3 U78 ( .A(n1), .Y(n74) );
  CLKINVX3 U79 ( .A(addr[6]), .Y(n75) );
endmodule


module crp_12 ( P, R, K_sub );
  output [1:32] P;
  input [1:32] R;
  input [1:48] K_sub;
  wire   n1;
  wire   [1:48] X;

  sbox1_12 u0 ( .addr(X[1:6]), .dout({P[9], P[17], P[23], P[31]}) );
  sbox2_12 u1 ( .addr({X[7], n1, X[9:12]}), .dout({P[13], P[28], P[2], P[18]})
         );
  sbox3_12 u2 ( .addr(X[13:18]), .dout({P[24], P[16], P[30], P[6]}) );
  sbox4_12 u3 ( .addr(X[19:24]), .dout({P[26], P[20], P[10], P[1]}) );
  sbox5_12 u4 ( .addr(X[25:30]), .dout({P[8], P[14], P[25], P[3]}) );
  sbox6_12 u5 ( .addr(X[31:36]), .dout({P[4], P[29], P[11], P[19]}) );
  sbox7_12 u6 ( .addr(X[37:42]), .dout({P[32], P[12], P[22], P[7]}) );
  sbox8_12 u7 ( .addr(X[43:48]), .dout({P[5], P[27], P[15], P[21]}) );
  XOR2X1 U1 ( .A(R[1]), .B(K_sub[2]), .Y(X[2]) );
  CLKXOR2X4 U2 ( .A(R[29]), .B(K_sub[42]), .Y(X[42]) );
  CLKXOR2X4 U3 ( .A(R[5]), .B(K_sub[6]), .Y(X[6]) );
  CLKXOR2X4 U4 ( .A(R[16]), .B(K_sub[25]), .Y(X[25]) );
  CLKXOR2X4 U5 ( .A(R[22]), .B(K_sub[33]), .Y(X[33]) );
  CLKXOR2X4 U6 ( .A(R[8]), .B(K_sub[11]), .Y(X[11]) );
  CLKXOR2X4 U7 ( .A(R[29]), .B(K_sub[44]), .Y(X[44]) );
  CLKXOR2X4 U8 ( .A(R[16]), .B(K_sub[23]), .Y(X[23]) );
  CLKXOR2X4 U9 ( .A(R[26]), .B(K_sub[39]), .Y(X[39]) );
  CLKXOR2X4 U10 ( .A(R[10]), .B(K_sub[15]), .Y(X[15]) );
  XNOR2X1 U11 ( .A(R[5]), .B(K_sub[8]), .Y(X[8]) );
  INVX3 U12 ( .A(X[8]), .Y(n1) );
  CLKXOR2X4 U13 ( .A(R[20]), .B(K_sub[31]), .Y(X[31]) );
  CLKXOR2X4 U14 ( .A(R[31]), .B(K_sub[46]), .Y(X[46]) );
  CLKXOR2X4 U15 ( .A(R[12]), .B(K_sub[19]), .Y(X[19]) );
  CLKXOR2X4 U16 ( .A(R[20]), .B(K_sub[29]), .Y(X[29]) );
  CLKXOR2X2 U17 ( .A(R[4]), .B(K_sub[5]), .Y(X[5]) );
  CLKXOR2X2 U18 ( .A(R[15]), .B(K_sub[22]), .Y(X[22]) );
  CLKXOR2X2 U19 ( .A(R[24]), .B(K_sub[35]), .Y(X[35]) );
  CLKXOR2X2 U20 ( .A(R[21]), .B(K_sub[30]), .Y(X[30]) );
  CLKXOR2X2 U21 ( .A(R[12]), .B(K_sub[17]), .Y(X[17]) );
  CLKXOR2X2 U22 ( .A(R[32]), .B(K_sub[1]), .Y(X[1]) );
  CLKXOR2X2 U23 ( .A(R[13]), .B(K_sub[20]), .Y(X[20]) );
  CLKXOR2X2 U24 ( .A(R[18]), .B(K_sub[27]), .Y(X[27]) );
  CLKXOR2X2 U25 ( .A(R[8]), .B(K_sub[13]), .Y(X[13]) );
  CLKXOR2X2 U26 ( .A(R[4]), .B(K_sub[7]), .Y(X[7]) );
  CLKXOR2X2 U27 ( .A(R[24]), .B(K_sub[37]), .Y(X[37]) );
  CLKXOR2X2 U28 ( .A(R[28]), .B(K_sub[43]), .Y(X[43]) );
  CLKXOR2X2 U29 ( .A(R[1]), .B(K_sub[48]), .Y(X[48]) );
  CLKXOR2X2 U30 ( .A(R[17]), .B(K_sub[24]), .Y(X[24]) );
  CLKXOR2X2 U31 ( .A(R[9]), .B(K_sub[12]), .Y(X[12]) );
  CLKXOR2X2 U32 ( .A(R[13]), .B(K_sub[18]), .Y(X[18]) );
  CLKXOR2X2 U33 ( .A(R[25]), .B(K_sub[36]), .Y(X[36]) );
  XOR2X1 U34 ( .A(R[23]), .B(K_sub[34]), .Y(X[34]) );
  XOR2X1 U35 ( .A(R[9]), .B(K_sub[14]), .Y(X[14]) );
  XOR2X1 U36 ( .A(R[30]), .B(K_sub[45]), .Y(X[45]) );
  XOR2X1 U37 ( .A(R[21]), .B(K_sub[32]), .Y(X[32]) );
  XOR2X1 U38 ( .A(R[25]), .B(K_sub[38]), .Y(X[38]) );
  XOR2X1 U39 ( .A(R[27]), .B(K_sub[40]), .Y(X[40]) );
  XOR2X1 U40 ( .A(R[3]), .B(K_sub[4]), .Y(X[4]) );
  XOR2X1 U41 ( .A(R[11]), .B(K_sub[16]), .Y(X[16]) );
  XOR2X1 U42 ( .A(R[7]), .B(K_sub[10]), .Y(X[10]) );
  XOR2X1 U43 ( .A(R[14]), .B(K_sub[21]), .Y(X[21]) );
  XOR2X1 U44 ( .A(R[6]), .B(K_sub[9]), .Y(X[9]) );
  XOR2X1 U45 ( .A(R[2]), .B(K_sub[3]), .Y(X[3]) );
  XOR2X1 U46 ( .A(R[28]), .B(K_sub[41]), .Y(X[41]) );
  XOR2X1 U47 ( .A(R[17]), .B(K_sub[26]), .Y(X[26]) );
  XOR2X1 U48 ( .A(R[32]), .B(K_sub[47]), .Y(X[47]) );
  XOR2X1 U49 ( .A(R[19]), .B(K_sub[28]), .Y(X[28]) );
endmodule


module sbox1_11 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127;

  OAI222X4 U13 ( .A0(addr[5]), .A1(n101), .B0(n1), .B1(n100), .C0(n99), .C1(n6), .Y(dout[3]) );
  OAI21X2 U42 ( .A0(n4), .A1(n112), .B0(n106), .Y(n123) );
  NAND2X2 U44 ( .A(addr[6]), .B(n10), .Y(n115) );
  NAND2X2 U48 ( .A(addr[1]), .B(n13), .Y(n114) );
  OAI22X2 U49 ( .A0(n69), .A1(n72), .B0(addr[5]), .B1(n120), .Y(n85) );
  NAND2X2 U50 ( .A(n3), .B(n69), .Y(n120) );
  NOR2X2 U51 ( .A(n69), .B(n3), .Y(n124) );
  NOR3X2 U55 ( .A(n2), .B(addr[6]), .C(n6), .Y(n102) );
  NOR2X2 U56 ( .A(n109), .B(n3), .Y(n93) );
  NAND2X2 U57 ( .A(addr[1]), .B(addr[6]), .Y(n109) );
  NAND2X2 U59 ( .A(n10), .B(n13), .Y(n112) );
  NOR2X1 U1 ( .A(n114), .B(n120), .Y(n104) );
  BUFX4 U2 ( .A(addr[4]), .Y(n2) );
  CLKBUFX3 U3 ( .A(addr[2]), .Y(n1) );
  OAI32X1 U4 ( .A0(n112), .A1(n2), .A2(n4), .B0(n115), .B1(n113), .Y(n80) );
  NOR2BXL U5 ( .AN(n118), .B(n1), .Y(n122) );
  CLKBUFX3 U6 ( .A(addr[2]), .Y(n4) );
  INVX3 U7 ( .A(addr[6]), .Y(n13) );
  OAI221X4 U8 ( .A0(addr[5]), .A1(n127), .B0(n126), .B1(n72), .C0(n125), .Y(
        dout[4]) );
  OAI221X4 U9 ( .A0(n88), .A1(n72), .B0(addr[5]), .B1(n87), .C0(n86), .Y(
        dout[2]) );
  OA21XL U10 ( .A0(n95), .A1(n115), .B0(n107), .Y(n119) );
  AOI222XL U11 ( .A0(n9), .A1(n1), .B0(n2), .B1(n110), .C0(n11), .C1(n6), .Y(
        n111) );
  AOI2BB2X1 U12 ( .B0(n2), .B1(n11), .A0N(addr[4]), .A1N(n115), .Y(n91) );
  BUFX4 U14 ( .A(addr[3]), .Y(n3) );
  CLKINVX1 U15 ( .A(n112), .Y(n9) );
  CLKINVX1 U16 ( .A(n113), .Y(n5) );
  NAND2BX1 U17 ( .AN(n104), .B(n119), .Y(n84) );
  CLKXOR2X2 U18 ( .A(n70), .B(n6), .Y(n90) );
  NOR2X1 U19 ( .A(n69), .B(n70), .Y(n118) );
  OAI21XL U20 ( .A0(n70), .A1(n114), .B0(n91), .Y(n92) );
  NAND2X1 U21 ( .A(n93), .B(n69), .Y(n107) );
  NAND2X1 U22 ( .A(n6), .B(n70), .Y(n113) );
  OAI211X1 U23 ( .A0(n69), .A1(n114), .B0(n108), .C0(n107), .Y(n89) );
  CLKINVX1 U24 ( .A(n109), .Y(n11) );
  NAND2X1 U25 ( .A(n124), .B(n8), .Y(n108) );
  CLKINVX1 U26 ( .A(n114), .Y(n12) );
  CLKINVX1 U27 ( .A(n115), .Y(n8) );
  CLKINVX1 U28 ( .A(n95), .Y(n71) );
  AO22X1 U29 ( .A0(n90), .A1(n8), .B0(n70), .B1(n123), .Y(n76) );
  OAI31X1 U30 ( .A0(n6), .A1(n3), .A2(n10), .B0(n103), .Y(n105) );
  AOI31XL U31 ( .A0(n10), .A1(n6), .A2(n2), .B0(n102), .Y(n103) );
  AOI211X1 U32 ( .A0(n7), .A1(n4), .B0(n117), .C0(n116), .Y(n126) );
  CLKINVX1 U33 ( .A(n108), .Y(n7) );
  AOI211X1 U34 ( .A0(n115), .A1(n114), .B0(n113), .C0(n2), .Y(n116) );
  OAI22X1 U35 ( .A0(n120), .A1(n112), .B0(n111), .B1(n70), .Y(n117) );
  AOI211X1 U36 ( .A0(n11), .A1(n118), .B0(n81), .C0(n80), .Y(n88) );
  OAI22X1 U37 ( .A0(n91), .A1(n6), .B0(n3), .B1(n106), .Y(n81) );
  CLKINVX3 U38 ( .A(addr[5]), .Y(n72) );
  NAND2X1 U39 ( .A(n3), .B(n72), .Y(n95) );
  NAND2X1 U40 ( .A(n12), .B(n1), .Y(n106) );
  XOR2X1 U41 ( .A(n82), .B(n2), .Y(n83) );
  NAND2X1 U43 ( .A(n1), .B(n3), .Y(n82) );
  OAI22XL U45 ( .A0(n3), .A1(n10), .B0(n70), .B1(n112), .Y(n94) );
  AOI211XL U46 ( .A0(n98), .A1(n70), .B0(n97), .C0(n104), .Y(n99) );
  OAI22XL U47 ( .A0(n96), .A1(n69), .B0(n95), .B1(n109), .Y(n97) );
  OAI22XL U52 ( .A0(n13), .A1(n72), .B0(n2), .B1(addr[1]), .Y(n98) );
  AOI221XL U53 ( .A0(n71), .A1(addr[6]), .B0(addr[5]), .B1(n94), .C0(n93), .Y(
        n96) );
  OAI21XL U54 ( .A0(addr[1]), .A1(n120), .B0(n119), .Y(n121) );
  AOI221XL U58 ( .A0(n9), .A1(n118), .B0(n93), .B1(n72), .C0(n75), .Y(n78) );
  OAI31X1 U60 ( .A0(n72), .A1(n2), .A2(n74), .B0(n73), .Y(n75) );
  OA21XL U61 ( .A0(n3), .A1(n13), .B0(n109), .Y(n74) );
  OAI21XL U62 ( .A0(n124), .A1(n85), .B0(n12), .Y(n73) );
  OAI21XL U63 ( .A0(n1), .A1(n10), .B0(n109), .Y(n110) );
  INVX4 U64 ( .A(n4), .Y(n6) );
  AOI222XL U65 ( .A0(n124), .A1(n123), .B0(n122), .B1(addr[6]), .C0(n1), .C1(
        n121), .Y(n125) );
  NOR4BBX1 U66 ( .AN(n107), .BN(n106), .C(n105), .D(n104), .Y(n127) );
  AOI222XL U67 ( .A0(n9), .A1(n90), .B0(n89), .B1(n6), .C0(n123), .C1(n69), 
        .Y(n101) );
  AOI2BB2XL U68 ( .B0(addr[5]), .B1(n92), .A0N(n120), .A1N(addr[1]), .Y(n100)
         );
  AOI32X1 U69 ( .A0(n4), .A1(n85), .A2(n9), .B0(n84), .B1(n6), .Y(n86) );
  AOI222XL U70 ( .A0(n124), .A1(n10), .B0(n83), .B1(addr[1]), .C0(n5), .C1(n13), .Y(n87) );
  OAI221X1 U71 ( .A0(n79), .A1(n72), .B0(n4), .B1(n78), .C0(n77), .Y(dout[1])
         );
  AOI32XL U72 ( .A0(addr[6]), .A1(n85), .A2(n1), .B0(n76), .B1(n72), .Y(n77)
         );
  AOI221X1 U73 ( .A0(n9), .A1(n90), .B0(n4), .B1(n93), .C0(n102), .Y(n79) );
  CLKINVX3 U74 ( .A(addr[1]), .Y(n10) );
  CLKINVX3 U75 ( .A(n2), .Y(n69) );
  CLKINVX3 U76 ( .A(n3), .Y(n70) );
endmodule


module sbox2_11 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147;

  NAND2X2 U55 ( .A(n2), .B(n8), .Y(n136) );
  NAND2X2 U57 ( .A(addr[2]), .B(n16), .Y(n104) );
  NAND2X2 U60 ( .A(addr[5]), .B(addr[2]), .Y(n132) );
  NOR2X2 U61 ( .A(n13), .B(n10), .Y(n101) );
  NAND2X2 U62 ( .A(n12), .B(n82), .Y(n146) );
  NAND2X2 U63 ( .A(n3), .B(n83), .Y(n124) );
  NAND2X2 U64 ( .A(addr[6]), .B(n12), .Y(n122) );
  NAND2X2 U67 ( .A(n3), .B(n2), .Y(n133) );
  AOI222XL U1 ( .A0(n4), .A1(n14), .B0(n88), .B1(n83), .C0(n140), .C1(n10), 
        .Y(n89) );
  CLKINVX1 U2 ( .A(n121), .Y(n13) );
  CLKINVX1 U3 ( .A(addr[5]), .Y(n1) );
  INVX3 U4 ( .A(addr[5]), .Y(n16) );
  OAI211X4 U5 ( .A0(n147), .A1(n146), .B0(n145), .C0(n144), .Y(dout[4]) );
  NAND3XL U6 ( .A(n98), .B(n97), .C(n96), .Y(dout[1]) );
  NAND2X1 U7 ( .A(addr[1]), .B(addr[6]), .Y(n121) );
  CLKINVX2 U8 ( .A(addr[1]), .Y(n12) );
  OAI221X1 U9 ( .A0(addr[1]), .A1(n136), .B0(n133), .B1(n12), .C0(n87), .Y(n95) );
  NOR2X1 U10 ( .A(n104), .B(n2), .Y(n141) );
  NOR2X1 U11 ( .A(n124), .B(n2), .Y(n140) );
  CLKBUFX4 U12 ( .A(addr[4]), .Y(n2) );
  NAND2X4 U13 ( .A(addr[1]), .B(n82), .Y(n114) );
  INVX3 U14 ( .A(addr[6]), .Y(n82) );
  NAND2XL U15 ( .A(n102), .B(n8), .Y(n109) );
  AOI211XL U16 ( .A0(n81), .A1(n95), .B0(n94), .C0(n93), .Y(n96) );
  AOI2BB2X1 U17 ( .B0(n16), .B1(n9), .A0N(n104), .A1N(n136), .Y(n117) );
  NOR3BXL U18 ( .AN(n135), .B(n134), .C(n4), .Y(n147) );
  BUFX4 U19 ( .A(addr[3]), .Y(n3) );
  NAND2X1 U20 ( .A(n4), .B(n13), .Y(n113) );
  CLKINVX1 U21 ( .A(n146), .Y(n10) );
  CLKINVX1 U22 ( .A(n115), .Y(n4) );
  CLKINVX1 U23 ( .A(n122), .Y(n11) );
  OAI31X1 U24 ( .A0(n124), .A1(n82), .A2(n16), .B0(n123), .Y(n128) );
  OAI21XL U25 ( .A0(n16), .A1(n12), .B0(n140), .Y(n123) );
  OAI22X1 U26 ( .A0(n122), .A1(n124), .B0(n101), .B1(n132), .Y(n84) );
  INVX1 U27 ( .A(n114), .Y(n14) );
  OAI22X1 U28 ( .A0(n122), .A1(n8), .B0(n5), .B1(n121), .Y(n129) );
  NAND3X1 U29 ( .A(n5), .B(n16), .C(n12), .Y(n111) );
  NAND2X1 U30 ( .A(n8), .B(n5), .Y(n115) );
  OAI21XL U31 ( .A0(n83), .A1(n133), .B0(n135), .Y(n85) );
  OAI22XL U32 ( .A0(n117), .A1(n146), .B0(n116), .B1(n132), .Y(n118) );
  AOI222XL U33 ( .A0(n14), .A1(n115), .B0(n6), .B1(n82), .C0(n4), .C1(n10), 
        .Y(n116) );
  CLKINVX1 U34 ( .A(n104), .Y(n15) );
  OAI2BB2XL U35 ( .B0(n114), .B1(n135), .A0N(n126), .A1N(n6), .Y(n106) );
  OAI21XL U36 ( .A0(n112), .A1(n114), .B0(n111), .Y(n120) );
  OAI21XL U37 ( .A0(n133), .A1(n114), .B0(n113), .Y(n119) );
  CLKINVX1 U38 ( .A(n124), .Y(n9) );
  CLKINVX1 U39 ( .A(n136), .Y(n7) );
  CLKINVX1 U40 ( .A(n133), .Y(n6) );
  CLKINVX1 U41 ( .A(n132), .Y(n81) );
  AOI2BB1X1 U42 ( .A0N(n126), .A1N(n125), .B0(n136), .Y(n127) );
  OAI22XL U43 ( .A0(n104), .A1(n114), .B0(n101), .B1(n132), .Y(n102) );
  AO21XL U44 ( .A0(n83), .A1(n7), .B0(n141), .Y(n86) );
  AO21X1 U45 ( .A0(n8), .A1(n15), .B0(n140), .Y(n142) );
  NAND3X1 U46 ( .A(n83), .B(n5), .C(addr[5]), .Y(n135) );
  OAI22X1 U47 ( .A0(addr[5]), .A1(n121), .B0(n122), .B1(n16), .Y(n126) );
  AOI2BB1X1 U48 ( .A0N(n3), .A1N(n1), .B0(n7), .Y(n112) );
  NOR3X1 U49 ( .A(addr[1]), .B(addr[2]), .C(n16), .Y(n125) );
  AOI2BB1XL U50 ( .A0N(n92), .A1N(n91), .B0(addr[5]), .Y(n93) );
  OAI22XL U51 ( .A0(n117), .A1(n114), .B0(n89), .B1(n1), .Y(n94) );
  OAI31XL U52 ( .A0(n114), .A1(n2), .A2(n8), .B0(n90), .Y(n91) );
  OAI21XL U53 ( .A0(n6), .A1(n9), .B0(n11), .Y(n90) );
  NAND2X1 U54 ( .A(n14), .B(n2), .Y(n137) );
  OAI31XL U56 ( .A0(n101), .A1(n3), .A2(addr[2]), .B0(n113), .Y(n92) );
  OAI211X1 U58 ( .A0(n139), .A1(n16), .B0(n138), .C0(n137), .Y(n143) );
  NAND3X1 U59 ( .A(n5), .B(n16), .C(addr[6]), .Y(n138) );
  AOI2BB2X1 U65 ( .B0(n11), .B1(n8), .A0N(n12), .A1N(n136), .Y(n139) );
  OAI22XL U66 ( .A0(addr[5]), .A1(n133), .B0(n3), .B1(n132), .Y(n134) );
  OAI2BB2XL U68 ( .B0(n112), .B1(n122), .A0N(n1), .A1N(n99), .Y(n100) );
  OAI211X1 U69 ( .A0(n146), .A1(n2), .B0(n137), .C0(n113), .Y(n99) );
  NAND3X1 U70 ( .A(n11), .B(n5), .C(n3), .Y(n87) );
  AOI2BB2XL U71 ( .B0(n3), .B1(n105), .A0N(n137), .A1N(n132), .Y(n108) );
  OAI211XL U72 ( .A0(n104), .A1(n146), .B0(n103), .C0(n111), .Y(n105) );
  NAND3XL U73 ( .A(addr[5]), .B(n5), .C(n13), .Y(n103) );
  OAI22XL U74 ( .A0(n3), .A1(n114), .B0(n82), .B1(n115), .Y(n88) );
  NAND4X1 U75 ( .A(n110), .B(n109), .C(n108), .D(n107), .Y(dout[2]) );
  AOI32XL U76 ( .A0(addr[1]), .A1(addr[2]), .A2(n7), .B0(n100), .B1(n83), .Y(
        n110) );
  AOI221XL U77 ( .A0(n125), .A1(addr[4]), .B0(n141), .B1(n11), .C0(n106), .Y(
        n107) );
  AOI33XL U78 ( .A0(n11), .A1(n15), .A2(n2), .B0(n81), .B1(n146), .B2(n3), .Y(
        n145) );
  AOI222XL U79 ( .A0(n143), .A1(n83), .B0(n13), .B1(n142), .C0(n14), .C1(n141), 
        .Y(n144) );
  AOI32XL U80 ( .A0(n15), .A1(n12), .A2(n4), .B0(n10), .B1(n86), .Y(n97) );
  AOI22X1 U81 ( .A0(n13), .A1(n85), .B0(n2), .B1(n84), .Y(n98) );
  NAND2X1 U82 ( .A(n131), .B(n130), .Y(dout[3]) );
  AOI221XL U83 ( .A0(n120), .A1(n83), .B0(addr[2]), .B1(n119), .C0(n118), .Y(
        n131) );
  AOI211X1 U84 ( .A0(n15), .A1(n129), .B0(n128), .C0(n127), .Y(n130) );
  CLKINVX3 U85 ( .A(n2), .Y(n5) );
  CLKINVX3 U86 ( .A(n3), .Y(n8) );
  CLKINVX3 U87 ( .A(addr[2]), .Y(n83) );
endmodule


module sbox3_11 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133;

  NOR2X2 U35 ( .A(n7), .B(addr[3]), .Y(n108) );
  NOR2X2 U50 ( .A(addr[1]), .B(addr[6]), .Y(n107) );
  NOR2X2 U52 ( .A(n76), .B(n2), .Y(n87) );
  NOR2X2 U56 ( .A(n76), .B(n78), .Y(n94) );
  NOR2X1 U1 ( .A(n7), .B(n76), .Y(n106) );
  OAI221X1 U2 ( .A0(n124), .A1(n7), .B0(n3), .B1(addr[1]), .C0(n19), .Y(n104)
         );
  OAI22XL U3 ( .A0(n2), .A1(n78), .B0(n3), .B1(n5), .Y(n123) );
  BUFX4 U4 ( .A(addr[4]), .Y(n2) );
  CLKBUFX3 U5 ( .A(n78), .Y(n1) );
  OAI33X1 U6 ( .A0(n9), .A1(n125), .A2(n78), .B0(n7), .B1(n94), .B2(n119), .Y(
        n79) );
  INVX3 U7 ( .A(n3), .Y(n78) );
  NOR2X1 U8 ( .A(n18), .B(n3), .Y(n91) );
  NOR2X1 U9 ( .A(n9), .B(n3), .Y(n121) );
  NOR2X1 U10 ( .A(n19), .B(n3), .Y(n95) );
  NOR2X1 U11 ( .A(n3), .B(n2), .Y(n110) );
  CLKBUFX4 U12 ( .A(addr[2]), .Y(n3) );
  OAI221X1 U13 ( .A0(addr[5]), .A1(n90), .B0(n89), .B1(n4), .C0(n88), .Y(
        dout[1]) );
  NOR2X4 U14 ( .A(n77), .B(n16), .Y(n124) );
  NOR2X4 U15 ( .A(addr[3]), .B(n2), .Y(n130) );
  NOR2X4 U16 ( .A(n16), .B(addr[6]), .Y(n125) );
  INVX3 U17 ( .A(addr[1]), .Y(n16) );
  NAND2XL U18 ( .A(n94), .B(n124), .Y(n132) );
  OAI211XL U19 ( .A0(n2), .A1(n17), .B0(n128), .C0(n127), .Y(n129) );
  NAND4XL U20 ( .A(n114), .B(n113), .C(n112), .D(n111), .Y(n115) );
  CLKINVX1 U21 ( .A(n132), .Y(n14) );
  INVX1 U22 ( .A(n124), .Y(n12) );
  CLKINVX1 U23 ( .A(n106), .Y(n5) );
  NAND2X1 U24 ( .A(n18), .B(n6), .Y(n122) );
  CLKINVX1 U25 ( .A(n86), .Y(n6) );
  CLKINVX1 U26 ( .A(n120), .Y(n20) );
  CLKINVX1 U27 ( .A(n119), .Y(n13) );
  CLKINVX1 U28 ( .A(n114), .Y(n10) );
  CLKINVX1 U29 ( .A(n107), .Y(n19) );
  NOR2X1 U30 ( .A(n18), .B(n78), .Y(n103) );
  NOR2X1 U31 ( .A(n12), .B(n78), .Y(n109) );
  INVX1 U32 ( .A(n125), .Y(n15) );
  AOI21X1 U33 ( .A0(n76), .A1(n78), .B0(n94), .Y(n120) );
  OAI21XL U34 ( .A0(n110), .A1(n130), .B0(n124), .Y(n82) );
  CLKINVX1 U36 ( .A(n81), .Y(n18) );
  NOR2X1 U37 ( .A(n15), .B(n7), .Y(n86) );
  NOR2X1 U38 ( .A(n124), .B(n107), .Y(n119) );
  OAI21XL U39 ( .A0(n109), .A1(n91), .B0(n130), .Y(n100) );
  NAND2X1 U40 ( .A(n103), .B(n87), .Y(n114) );
  CLKINVX1 U41 ( .A(n87), .Y(n9) );
  CLKINVX1 U42 ( .A(n91), .Y(n17) );
  CLKINVX1 U43 ( .A(n110), .Y(n11) );
  CLKINVX1 U44 ( .A(n121), .Y(n8) );
  OR2X1 U45 ( .A(n103), .B(n95), .Y(n126) );
  OAI221X1 U46 ( .A0(n15), .A1(n11), .B0(n78), .B1(n6), .C0(n93), .Y(n98) );
  AOI221XL U47 ( .A0(n95), .A1(n2), .B0(n92), .B1(n7), .C0(n14), .Y(n93) );
  OAI21XL U48 ( .A0(n1), .A1(n19), .B0(n17), .Y(n92) );
  XNOR2X1 U49 ( .A(addr[5]), .B(addr[3]), .Y(n102) );
  CLKINVX1 U51 ( .A(addr[5]), .Y(n4) );
  OAI221X1 U53 ( .A0(n19), .A1(n11), .B0(n12), .B1(n9), .C0(n105), .Y(n116) );
  AOI221XL U54 ( .A0(addr[3]), .A1(n104), .B0(n103), .B1(n130), .C0(n14), .Y(
        n105) );
  CLKINVX1 U55 ( .A(addr[6]), .Y(n77) );
  NAND3X1 U57 ( .A(n3), .B(n16), .C(n108), .Y(n113) );
  NOR2X1 U58 ( .A(n77), .B(addr[1]), .Y(n81) );
  AOI32XL U59 ( .A0(n1), .A1(n76), .A2(n124), .B0(n123), .B1(n77), .Y(n128) );
  AOI22XL U60 ( .A0(n2), .A1(n126), .B0(n125), .B1(n130), .Y(n127) );
  AOI222XL U61 ( .A0(n110), .A1(n125), .B0(n109), .B1(n76), .C0(n108), .C1(
        n107), .Y(n111) );
  OAI211XL U62 ( .A0(n106), .A1(n130), .B0(n1), .C0(addr[6]), .Y(n112) );
  OAI21XL U63 ( .A0(n3), .A1(addr[1]), .B0(n15), .Y(n80) );
  AOI221XL U64 ( .A0(n86), .A1(n76), .B0(n87), .B1(n125), .C0(n85), .Y(n89) );
  OAI211X1 U65 ( .A0(n84), .A1(n78), .B0(n83), .C0(n82), .Y(n85) );
  AOI222XL U66 ( .A0(n81), .A1(n76), .B0(n107), .B1(n106), .C0(n130), .C1(n16), 
        .Y(n84) );
  OAI21XL U67 ( .A0(n91), .A1(n14), .B0(addr[4]), .Y(n83) );
  AOI221XL U68 ( .A0(n125), .A1(n20), .B0(addr[3]), .B1(n126), .C0(n96), .Y(
        n97) );
  OAI22X1 U69 ( .A0(n12), .A1(n8), .B0(n5), .B1(n18), .Y(n96) );
  OAI211X1 U70 ( .A0(n19), .A1(n8), .B0(n118), .C0(n117), .Y(dout[3]) );
  AOI32XL U71 ( .A0(n125), .A1(n3), .A2(n102), .B0(n108), .B1(n109), .Y(n118)
         );
  AOI22XL U72 ( .A0(n116), .A1(n4), .B0(addr[5]), .B1(n115), .Y(n117) );
  AOI221XL U73 ( .A0(n121), .A1(n125), .B0(n95), .B1(n108), .C0(n10), .Y(n88)
         );
  AOI221XL U74 ( .A0(n130), .A1(n80), .B0(n94), .B1(n122), .C0(n79), .Y(n90)
         );
  NAND4X1 U75 ( .A(n101), .B(n113), .C(n100), .D(n99), .Y(dout[2]) );
  NAND3XL U76 ( .A(n2), .B(n124), .C(n102), .Y(n101) );
  AOI2BB2XL U77 ( .B0(addr[5]), .B1(n98), .A0N(addr[5]), .A1N(n97), .Y(n99) );
  OAI221X1 U78 ( .A0(n133), .A1(n4), .B0(n2), .B1(n132), .C0(n131), .Y(dout[4]) );
  AOI32XL U79 ( .A0(n130), .A1(n77), .A2(addr[2]), .B0(n129), .B1(n4), .Y(n131) );
  AOI222XL U80 ( .A0(n20), .A1(n122), .B0(n121), .B1(addr[1]), .C0(n120), .C1(
        n13), .Y(n133) );
  CLKINVX3 U81 ( .A(n2), .Y(n7) );
  CLKINVX3 U82 ( .A(addr[3]), .Y(n76) );
endmodule


module sbox4_11 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126;

  OAI32X4 U12 ( .A0(n12), .A1(n2), .A2(addr[2]), .B0(n11), .B1(n108), .Y(n123)
         );
  OAI222X4 U20 ( .A0(addr[2]), .A1(n92), .B0(n106), .B1(n91), .C0(n90), .C1(
        n72), .Y(dout[2]) );
  OAI222X4 U33 ( .A0(addr[4]), .A1(n106), .B0(n6), .B1(n108), .C0(n2), .C1(
        n118), .Y(n83) );
  NAND2X2 U34 ( .A(addr[4]), .B(n2), .Y(n108) );
  NOR2X2 U43 ( .A(n71), .B(addr[4]), .Y(n113) );
  NOR2X2 U45 ( .A(n11), .B(n2), .Y(n111) );
  NAND2X2 U51 ( .A(n6), .B(n14), .Y(n118) );
  NOR2X2 U52 ( .A(n16), .B(addr[5]), .Y(n97) );
  NAND2X2 U53 ( .A(addr[6]), .B(addr[1]), .Y(n85) );
  NAND2X2 U54 ( .A(addr[1]), .B(n14), .Y(n116) );
  NOR2X2 U55 ( .A(n115), .B(n11), .Y(n121) );
  NAND2X2 U56 ( .A(n71), .B(n16), .Y(n115) );
  NAND2X2 U57 ( .A(addr[5]), .B(n16), .Y(n96) );
  NAND2X2 U58 ( .A(addr[6]), .B(n6), .Y(n106) );
  OAI222X1 U1 ( .A0(n12), .A1(n85), .B0(n97), .B1(n116), .C0(n16), .C1(n118), 
        .Y(n73) );
  CLKINVX1 U2 ( .A(n116), .Y(n9) );
  OAI31X4 U3 ( .A0(n118), .A1(n11), .A2(n16), .B0(n117), .Y(n119) );
  CLKINVX1 U4 ( .A(n71), .Y(n1) );
  CLKBUFX3 U5 ( .A(addr[3]), .Y(n2) );
  OAI221X1 U6 ( .A0(addr[2]), .A1(n80), .B0(n118), .B1(n105), .C0(n79), .Y(
        dout[1]) );
  INVX4 U7 ( .A(addr[5]), .Y(n11) );
  OAI31X1 U8 ( .A0(n108), .A1(addr[5]), .A2(n5), .B0(n107), .Y(n109) );
  AOI222XL U9 ( .A0(n16), .A1(n14), .B0(n113), .B1(n6), .C0(addr[1]), .C1(n71), 
        .Y(n114) );
  OAI222X1 U10 ( .A0(addr[1]), .A1(n84), .B0(n85), .B1(n74), .C0(n71), .C1(
        n107), .Y(n75) );
  NAND2XL U11 ( .A(n1), .B(addr[5]), .Y(n84) );
  AOI211XL U13 ( .A0(n83), .A1(n11), .B0(n82), .C0(n7), .Y(n92) );
  NAND2XL U14 ( .A(n16), .B(n11), .Y(n74) );
  CLKINVX1 U15 ( .A(n118), .Y(n3) );
  CLKINVX1 U16 ( .A(n115), .Y(n15) );
  CLKINVX1 U17 ( .A(n112), .Y(n4) );
  OAI21X1 U18 ( .A0(n9), .A1(n5), .B0(n72), .Y(n112) );
  AOI22X1 U19 ( .A0(n10), .A1(n111), .B0(n5), .B1(n113), .Y(n93) );
  OAI211X1 U21 ( .A0(n6), .A1(n115), .B0(n93), .C0(n8), .Y(n94) );
  CLKINVX1 U22 ( .A(n85), .Y(n10) );
  NAND2X1 U23 ( .A(n97), .B(n71), .Y(n105) );
  NAND2X1 U24 ( .A(n113), .B(n3), .Y(n98) );
  NAND2X1 U25 ( .A(n9), .B(n97), .Y(n107) );
  NAND2X1 U26 ( .A(n118), .B(n85), .Y(n110) );
  OAI21XL U27 ( .A0(n15), .A1(n11), .B0(n108), .Y(n95) );
  CLKINVX1 U28 ( .A(n84), .Y(n13) );
  CLKINVX1 U29 ( .A(addr[2]), .Y(n72) );
  OAI31X1 U30 ( .A0(n16), .A1(addr[6]), .A2(n11), .B0(n87), .Y(n88) );
  OAI21XL U31 ( .A0(n113), .A1(n12), .B0(n10), .Y(n87) );
  OAI211X1 U32 ( .A0(n76), .A1(n16), .B0(n98), .C0(n8), .Y(n77) );
  AOI222XL U35 ( .A0(addr[5]), .A1(addr[6]), .B0(n111), .B1(addr[1]), .C0(n5), 
        .C1(n2), .Y(n76) );
  NAND3XL U36 ( .A(n10), .B(n71), .C(addr[4]), .Y(n117) );
  OAI22XL U37 ( .A0(n116), .A1(n115), .B0(n1), .B1(n112), .Y(n78) );
  CLKINVX3 U38 ( .A(addr[4]), .Y(n16) );
  OAI2BB2XL U39 ( .B0(n115), .B1(n106), .A0N(n11), .A1N(n86), .Y(n89) );
  OAI221XL U40 ( .A0(n116), .A1(addr[4]), .B0(n108), .B1(addr[1]), .C0(n117), 
        .Y(n86) );
  CLKINVX1 U41 ( .A(addr[6]), .Y(n14) );
  CLKINVX1 U42 ( .A(n81), .Y(n7) );
  OAI21XL U44 ( .A0(n96), .A1(n118), .B0(n93), .Y(n82) );
  NAND3X1 U46 ( .A(n101), .B(n100), .C(n99), .Y(n102) );
  AOI32X1 U47 ( .A0(n96), .A1(n71), .A2(n9), .B0(n10), .B1(n95), .Y(n101) );
  AOI2BB2XL U48 ( .B0(n6), .B1(n121), .A0N(n98), .A1N(addr[5]), .Y(n99) );
  OAI21XL U49 ( .A0(n97), .A1(n12), .B0(n5), .Y(n100) );
  AOI2BB2XL U50 ( .B0(n5), .B1(n123), .A0N(n122), .A1N(n72), .Y(n124) );
  AOI211XL U59 ( .A0(n5), .A1(n121), .B0(n120), .C0(n119), .Y(n122) );
  OAI22XL U60 ( .A0(n116), .A1(n115), .B0(addr[5]), .B1(n114), .Y(n120) );
  CLKINVX1 U61 ( .A(n75), .Y(n8) );
  AOI32XL U62 ( .A0(n9), .A1(n96), .A2(n1), .B0(addr[1]), .B1(n121), .Y(n81)
         );
  AOI222XL U63 ( .A0(n5), .A1(n12), .B0(n121), .B1(n116), .C0(n2), .C1(n73), 
        .Y(n80) );
  AOI22XL U64 ( .A0(n78), .A1(n11), .B0(addr[2]), .B1(n77), .Y(n79) );
  NAND2XL U65 ( .A(n111), .B(addr[4]), .Y(n91) );
  AOI211X1 U66 ( .A0(n13), .A1(n110), .B0(n89), .C0(n88), .Y(n90) );
  OAI211X1 U67 ( .A0(n106), .A1(n105), .B0(n104), .C0(n103), .Y(dout[3]) );
  AOI32X1 U68 ( .A0(n2), .A1(n12), .A2(n9), .B0(n94), .B1(n72), .Y(n104) );
  AOI22XL U69 ( .A0(addr[2]), .A1(n102), .B0(n3), .B1(n123), .Y(n103) );
  OAI211X1 U70 ( .A0(addr[2]), .A1(n126), .B0(n125), .C0(n124), .Y(dout[4]) );
  AOI32X1 U71 ( .A0(n10), .A1(n12), .A2(n2), .B0(n4), .B1(n13), .Y(n125) );
  AOI221XL U72 ( .A0(n3), .A1(n111), .B0(n15), .B1(n110), .C0(n109), .Y(n126)
         );
  CLKINVX3 U73 ( .A(n106), .Y(n5) );
  CLKINVX3 U74 ( .A(addr[1]), .Y(n6) );
  CLKINVX3 U75 ( .A(n96), .Y(n12) );
  CLKINVX3 U76 ( .A(n2), .Y(n71) );
endmodule


module sbox5_11 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121;

  OAI222X4 U18 ( .A0(addr[3]), .A1(n106), .B0(n69), .B1(n90), .C0(n14), .C1(n9), .Y(n93) );
  OAI22X2 U40 ( .A0(addr[5]), .A1(n106), .B0(n70), .B1(n114), .Y(n116) );
  NOR2X2 U41 ( .A(n3), .B(addr[3]), .Y(n102) );
  NAND2X2 U45 ( .A(addr[6]), .B(n9), .Y(n114) );
  NAND2X2 U50 ( .A(n9), .B(n69), .Y(n110) );
  NAND2X2 U52 ( .A(addr[1]), .B(n69), .Y(n113) );
  NAND2X2 U54 ( .A(addr[1]), .B(addr[6]), .Y(n106) );
  NAND2X2 U55 ( .A(addr[3]), .B(n14), .Y(n121) );
  CLKINVX1 U1 ( .A(addr[5]), .Y(n1) );
  AOI221XL U2 ( .A0(n93), .A1(n1), .B0(n10), .B1(n15), .C0(n92), .Y(n105) );
  INVX3 U3 ( .A(addr[5]), .Y(n70) );
  OAI221X4 U4 ( .A0(n111), .A1(n110), .B0(n121), .B1(n114), .C0(n109), .Y(n112) );
  OAI221X4 U5 ( .A0(n14), .A1(n114), .B0(n70), .B1(n113), .C0(n120), .Y(n115)
         );
  OAI221X4 U6 ( .A0(n107), .A1(n121), .B0(n111), .B1(n113), .C0(n85), .Y(n86)
         );
  OAI31X1 U7 ( .A0(n68), .A1(addr[5]), .A2(addr[1]), .B0(n81), .Y(n73) );
  OAI32X1 U8 ( .A0(n114), .A1(addr[5]), .A2(n3), .B0(n13), .B1(n107), .Y(n79)
         );
  AOI32XL U9 ( .A0(n15), .A1(n98), .A2(n12), .B0(n2), .B1(n73), .Y(n77) );
  CLKBUFX3 U10 ( .A(addr[4]), .Y(n2) );
  CLKINVX1 U11 ( .A(n81), .Y(n5) );
  NAND2X1 U12 ( .A(n6), .B(n15), .Y(n81) );
  CLKINVX1 U13 ( .A(n110), .Y(n8) );
  CLKXOR2X2 U14 ( .A(n68), .B(n70), .Y(n94) );
  AOI2BB1X1 U15 ( .A0N(n14), .A1N(n1), .B0(n15), .Y(n111) );
  NOR2X1 U16 ( .A(n121), .B(n70), .Y(n91) );
  NOR2BX1 U17 ( .AN(n116), .B(n90), .Y(n83) );
  NAND2X1 U19 ( .A(n8), .B(n70), .Y(n120) );
  CLKINVX1 U20 ( .A(n113), .Y(n12) );
  NAND2X1 U21 ( .A(n12), .B(n70), .Y(n107) );
  CLKINVX1 U22 ( .A(n121), .Y(n13) );
  OAI31X1 U23 ( .A0(n4), .A1(n15), .A2(n113), .B0(n99), .Y(n72) );
  CLKINVX1 U24 ( .A(n106), .Y(n10) );
  OAI2BB2XL U25 ( .B0(n1), .B1(n113), .A0N(n98), .A1N(n6), .Y(n101) );
  CLKINVX1 U26 ( .A(n114), .Y(n6) );
  CLKINVX1 U27 ( .A(n90), .Y(n16) );
  CLKINVX1 U28 ( .A(addr[1]), .Y(n9) );
  CLKINVX1 U29 ( .A(addr[3]), .Y(n68) );
  CLKINVX1 U30 ( .A(addr[6]), .Y(n69) );
  AOI211X1 U31 ( .A0(n91), .A1(addr[1]), .B0(n80), .C0(n79), .Y(n89) );
  OAI2BB2XL U32 ( .B0(n111), .B1(n106), .A0N(n94), .A1N(n8), .Y(n80) );
  AOI211X1 U33 ( .A0(n102), .A1(n84), .B0(n83), .C0(n82), .Y(n85) );
  OAI21XL U34 ( .A0(n69), .A1(n1), .B0(n106), .Y(n84) );
  NOR3XL U35 ( .A(n94), .B(n3), .C(n110), .Y(n82) );
  AOI222XL U36 ( .A0(n10), .A1(n16), .B0(addr[5]), .B1(n108), .C0(n11), .C1(
        n14), .Y(n109) );
  CLKINVX1 U37 ( .A(n107), .Y(n11) );
  OAI21XL U38 ( .A0(addr[6]), .A1(addr[3]), .B0(n106), .Y(n108) );
  NAND2X1 U39 ( .A(addr[3]), .B(n3), .Y(n90) );
  NAND2X1 U42 ( .A(n2), .B(addr[5]), .Y(n98) );
  NAND2X1 U43 ( .A(n3), .B(n68), .Y(n97) );
  OAI21XL U44 ( .A0(addr[1]), .A1(n97), .B0(n96), .Y(n103) );
  AOI33XL U46 ( .A0(n3), .A1(n95), .A2(addr[5]), .B0(n94), .B1(n14), .B2(
        addr[1]), .Y(n96) );
  OAI21XL U47 ( .A0(n9), .A1(n68), .B0(n114), .Y(n95) );
  OAI21XL U48 ( .A0(addr[6]), .A1(n121), .B0(n99), .Y(n100) );
  NAND2X1 U49 ( .A(n71), .B(n8), .Y(n99) );
  XOR2X1 U51 ( .A(n4), .B(n3), .Y(n71) );
  AOI2BB2XL U53 ( .B0(n102), .B1(n116), .A0N(n2), .A1N(n75), .Y(n76) );
  AOI211X1 U56 ( .A0(n7), .A1(n3), .B0(n74), .C0(n83), .Y(n75) );
  AO22XL U57 ( .A0(n12), .A1(n13), .B0(addr[6]), .B1(n102), .Y(n74) );
  CLKINVX1 U58 ( .A(n120), .Y(n7) );
  CLKINVX1 U59 ( .A(n2), .Y(n4) );
  AO22XL U60 ( .A0(n12), .A1(n16), .B0(addr[6]), .B1(n91), .Y(n92) );
  AOI222XL U61 ( .A0(n116), .A1(n14), .B0(addr[3]), .B1(n115), .C0(n12), .C1(
        n15), .Y(n117) );
  OAI221X1 U62 ( .A0(n2), .A1(n105), .B0(n110), .B1(n121), .C0(n104), .Y(
        dout[3]) );
  AOI222XL U63 ( .A0(n2), .A1(n103), .B0(n102), .B1(n101), .C0(n100), .C1(n1), 
        .Y(n104) );
  OAI211X1 U64 ( .A0(n2), .A1(n89), .B0(n88), .C0(n87), .Y(dout[2]) );
  AOI33XL U65 ( .A0(n13), .A1(n98), .A2(n6), .B0(n3), .B1(n94), .B2(n8), .Y(
        n88) );
  AOI222XL U66 ( .A0(n5), .A1(n70), .B0(n2), .B1(n86), .C0(n91), .C1(n10), .Y(
        n87) );
  OAI211X1 U67 ( .A0(n78), .A1(n70), .B0(n77), .C0(n76), .Y(dout[1]) );
  AOI221XL U68 ( .A0(n13), .A1(addr[1]), .B0(n10), .B1(n15), .C0(n72), .Y(n78)
         );
  OAI211X1 U69 ( .A0(n121), .A1(n120), .B0(n119), .C0(n118), .Y(dout[4]) );
  AOI32XL U70 ( .A0(n15), .A1(n114), .A2(addr[5]), .B0(n2), .B1(n112), .Y(n119) );
  AOI2BB2X1 U71 ( .B0(n5), .B1(n70), .A0N(n2), .A1N(n117), .Y(n118) );
  BUFX4 U72 ( .A(addr[2]), .Y(n3) );
  CLKINVX3 U73 ( .A(n3), .Y(n14) );
  CLKINVX3 U74 ( .A(n97), .Y(n15) );
endmodule


module sbox6_11 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147;

  NAND2X2 U39 ( .A(n138), .B(addr[3]), .Y(n147) );
  NOR2X2 U47 ( .A(n15), .B(n81), .Y(n138) );
  NOR2X2 U50 ( .A(n17), .B(n4), .Y(n119) );
  NOR2X2 U58 ( .A(n11), .B(n17), .Y(n125) );
  NAND2X2 U61 ( .A(n97), .B(n103), .Y(n112) );
  NOR2X2 U62 ( .A(n85), .B(addr[1]), .Y(n103) );
  NOR2X2 U63 ( .A(n11), .B(addr[3]), .Y(n97) );
  NAND2X2 U64 ( .A(n117), .B(n131), .Y(n140) );
  NOR2X2 U65 ( .A(n5), .B(addr[3]), .Y(n131) );
  NOR2X2 U66 ( .A(n82), .B(addr[6]), .Y(n117) );
  NOR2X1 U1 ( .A(n15), .B(addr[3]), .Y(n102) );
  AOI211X1 U2 ( .A0(n7), .A1(n17), .B0(n131), .C0(n143), .Y(n121) );
  CLKINVX1 U3 ( .A(addr[3]), .Y(n1) );
  INVX3 U4 ( .A(addr[3]), .Y(n17) );
  CLKINVX1 U5 ( .A(n15), .Y(n2) );
  OAI222X1 U6 ( .A0(n91), .A1(n7), .B0(n5), .B1(n10), .C0(addr[5]), .C1(n12), 
        .Y(n92) );
  BUFX4 U7 ( .A(addr[2]), .Y(n5) );
  CLKINVX1 U8 ( .A(n11), .Y(n3) );
  INVX4 U9 ( .A(n4), .Y(n11) );
  CLKBUFX3 U10 ( .A(addr[4]), .Y(n4) );
  OAI221X1 U11 ( .A0(n85), .A1(n9), .B0(n17), .B1(n18), .C0(n86), .Y(n90) );
  INVX3 U12 ( .A(n96), .Y(n18) );
  OAI221X4 U13 ( .A0(n123), .A1(n83), .B0(n81), .B1(n7), .C0(n16), .Y(n124) );
  NOR2X4 U14 ( .A(addr[1]), .B(addr[6]), .Y(n130) );
  NOR2X4 U15 ( .A(n5), .B(addr[5]), .Y(n143) );
  INVX1 U16 ( .A(n130), .Y(n84) );
  CLKINVX1 U17 ( .A(n125), .Y(n9) );
  NAND2X1 U18 ( .A(n84), .B(n18), .Y(n105) );
  INVXL U19 ( .A(n121), .Y(n6) );
  CLKINVX1 U20 ( .A(n138), .Y(n14) );
  CLKINVX1 U21 ( .A(n117), .Y(n81) );
  CLKINVX1 U22 ( .A(n119), .Y(n12) );
  NOR2X1 U23 ( .A(n18), .B(n123), .Y(n144) );
  NOR2X1 U24 ( .A(n82), .B(n85), .Y(n96) );
  CLKINVX1 U25 ( .A(n103), .Y(n83) );
  OAI211X1 U26 ( .A0(n84), .A1(n9), .B0(n104), .C0(n112), .Y(n108) );
  OAI21XL U27 ( .A0(n103), .A1(n117), .B0(n102), .Y(n104) );
  OAI21XL U28 ( .A0(n132), .A1(n85), .B0(n1), .Y(n86) );
  AOI21X1 U29 ( .A0(n11), .A1(n102), .B0(n125), .Y(n91) );
  OAI2BB2XL U30 ( .B0(n143), .B1(n84), .A0N(n143), .A1N(n117), .Y(n118) );
  CLKINVX1 U31 ( .A(n122), .Y(n16) );
  CLKINVX1 U32 ( .A(n126), .Y(n13) );
  CLKINVX1 U33 ( .A(n97), .Y(n10) );
  NAND2BX1 U34 ( .AN(n144), .B(n137), .Y(n107) );
  CLKINVX1 U35 ( .A(addr[1]), .Y(n82) );
  NOR2X1 U36 ( .A(n18), .B(n2), .Y(n122) );
  NOR2X1 U37 ( .A(addr[1]), .B(n3), .Y(n132) );
  OAI22X1 U38 ( .A0(n12), .A1(n81), .B0(n5), .B1(n13), .Y(n88) );
  NAND2X1 U40 ( .A(n2), .B(n7), .Y(n123) );
  NAND4X1 U41 ( .A(n147), .B(n140), .C(n100), .D(n99), .Y(n101) );
  AOI222XL U42 ( .A0(n98), .A1(n15), .B0(n102), .B1(n130), .C0(n97), .C1(n105), 
        .Y(n99) );
  NAND3X1 U43 ( .A(n5), .B(n12), .C(n96), .Y(n100) );
  OAI221X1 U44 ( .A0(n17), .A1(n83), .B0(n12), .B1(n85), .C0(n13), .Y(n98) );
  AOI22X1 U45 ( .A0(n4), .A1(n115), .B0(addr[5]), .B1(n114), .Y(n129) );
  OAI21XL U46 ( .A0(n121), .A1(n84), .B0(n147), .Y(n115) );
  OAI21XL U48 ( .A0(n113), .A1(n15), .B0(n112), .Y(n114) );
  AOI221XL U49 ( .A0(n119), .A1(n82), .B0(n130), .B1(addr[3]), .C0(n111), .Y(
        n113) );
  OAI22XL U51 ( .A0(n81), .A1(n11), .B0(addr[3]), .B1(n18), .Y(n111) );
  OAI22XL U52 ( .A0(n17), .A1(n85), .B0(addr[1]), .B1(n12), .Y(n142) );
  AOI211X1 U53 ( .A0(n4), .A1(n135), .B0(n134), .C0(n133), .Y(n136) );
  OA21XL U54 ( .A0(n1), .A1(n2), .B0(n132), .Y(n133) );
  OAI2BB2XL U55 ( .B0(n3), .B1(n16), .A0N(n131), .A1N(n130), .Y(n134) );
  OAI22X1 U56 ( .A0(n5), .A1(n81), .B0(n15), .B1(n18), .Y(n135) );
  CLKINVX3 U57 ( .A(addr[5]), .Y(n7) );
  AOI2BB2X1 U59 ( .B0(n5), .B1(n130), .A0N(n2), .A1N(n83), .Y(n137) );
  NOR2X1 U60 ( .A(n83), .B(n3), .Y(n126) );
  AOI2BB2XL U67 ( .B0(n143), .B1(n90), .A0N(n89), .A1N(n7), .Y(n94) );
  AOI211X1 U68 ( .A0(n122), .A1(n4), .B0(n88), .C0(n87), .Y(n89) );
  OAI32X1 U69 ( .A0(n83), .A1(n17), .A2(n15), .B0(n14), .B1(n10), .Y(n87) );
  NAND3X1 U70 ( .A(n147), .B(n140), .C(n139), .Y(n141) );
  AOI32X1 U71 ( .A0(n5), .A1(n82), .A2(n4), .B0(n138), .B1(n11), .Y(n139) );
  AO22XL U72 ( .A0(n143), .A1(n3), .B0(n116), .B1(n11), .Y(n120) );
  OAI21XL U73 ( .A0(n2), .A1(n7), .B0(n123), .Y(n116) );
  CLKINVX1 U74 ( .A(n106), .Y(n8) );
  AOI32XL U75 ( .A0(n105), .A1(n11), .A2(n1), .B0(addr[1]), .B1(n125), .Y(n106) );
  OAI211X1 U76 ( .A0(n11), .A1(n140), .B0(n110), .C0(n109), .Y(dout[2]) );
  AOI222XL U77 ( .A0(n108), .A1(n7), .B0(n143), .B1(n8), .C0(n119), .C1(n107), 
        .Y(n109) );
  AOI2BB2XL U78 ( .B0(addr[5]), .B1(n101), .A0N(n15), .A1N(n112), .Y(n110) );
  OAI211X1 U79 ( .A0(n3), .A1(n147), .B0(n146), .C0(n145), .Y(dout[4]) );
  AOI222XL U80 ( .A0(n144), .A1(n17), .B0(n143), .B1(n142), .C0(n141), .C1(n7), 
        .Y(n145) );
  OA22X1 U81 ( .A0(n9), .A1(n137), .B0(n136), .B1(n7), .Y(n146) );
  NAND3X1 U82 ( .A(n129), .B(n128), .C(n127), .Y(dout[3]) );
  AOI32XL U83 ( .A0(n120), .A1(n17), .A2(addr[1]), .B0(n119), .B1(n118), .Y(
        n128) );
  AOI222XL U84 ( .A0(n144), .A1(n11), .B0(n126), .B1(n6), .C0(n125), .C1(n124), 
        .Y(n127) );
  NAND3BX1 U85 ( .AN(n95), .B(n94), .C(n93), .Y(dout[1]) );
  OAI222X1 U86 ( .A0(n140), .A1(n4), .B0(n112), .B1(n15), .C0(n18), .C1(n91), 
        .Y(n95) );
  AOI32XL U87 ( .A0(addr[1]), .A1(n7), .A2(n125), .B0(n130), .B1(n92), .Y(n93)
         );
  CLKINVX3 U88 ( .A(n5), .Y(n15) );
  CLKINVX3 U89 ( .A(addr[6]), .Y(n85) );
endmodule


module sbox7_11 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148;

  OAI222X4 U19 ( .A0(n20), .A1(n129), .B0(n4), .B1(n17), .C0(addr[1]), .C1(n85), .Y(n122) );
  OAI33X4 U33 ( .A0(addr[1]), .A1(n4), .A2(n5), .B0(n18), .B1(n86), .B2(n83), 
        .Y(n97) );
  NOR2X2 U44 ( .A(n84), .B(n4), .Y(n116) );
  NOR2X2 U48 ( .A(addr[1]), .B(addr[6]), .Y(n136) );
  NOR2X2 U51 ( .A(n10), .B(n84), .Y(n125) );
  NOR2X2 U52 ( .A(n18), .B(addr[3]), .Y(n131) );
  NOR2X2 U58 ( .A(n93), .B(n124), .Y(n142) );
  NOR2X2 U60 ( .A(n19), .B(addr[1]), .Y(n93) );
  NOR2X2 U62 ( .A(n87), .B(n3), .Y(n137) );
  NOR2X2 U65 ( .A(n19), .B(n21), .Y(n140) );
  NAND2X1 U1 ( .A(n3), .B(n4), .Y(n119) );
  CLKBUFX3 U2 ( .A(addr[4]), .Y(n4) );
  CLKINVX1 U3 ( .A(n87), .Y(n1) );
  CLKINVX1 U4 ( .A(n86), .Y(n2) );
  CLKBUFX3 U5 ( .A(addr[2]), .Y(n5) );
  OAI31X1 U6 ( .A0(n84), .A1(n87), .A2(n21), .B0(n117), .Y(n121) );
  NOR2X4 U7 ( .A(n21), .B(addr[6]), .Y(n124) );
  OAI22X1 U8 ( .A0(addr[1]), .A1(n85), .B0(n5), .B1(n113), .Y(n100) );
  OAI22X1 U9 ( .A0(n4), .A1(n10), .B0(addr[3]), .B1(n13), .Y(n103) );
  AOI211XL U10 ( .A0(n5), .A1(n16), .B0(n131), .C0(n130), .Y(n132) );
  NOR3XL U11 ( .A(n20), .B(addr[3]), .C(n2), .Y(n130) );
  OAI21XL U12 ( .A0(n3), .A1(n1), .B0(n119), .Y(n89) );
  BUFX4 U13 ( .A(addr[5]), .Y(n3) );
  AOI221XL U14 ( .A0(n140), .A1(n89), .B0(n109), .B1(n16), .C0(n88), .Y(n96)
         );
  CLKINVX1 U15 ( .A(n140), .Y(n18) );
  OAI2BB2XL U16 ( .B0(n142), .B1(n13), .A0N(n141), .A1N(n140), .Y(n143) );
  CLKINVX1 U17 ( .A(n125), .Y(n8) );
  CLKINVX1 U18 ( .A(n142), .Y(n16) );
  NAND2X1 U20 ( .A(n8), .B(n14), .Y(n105) );
  CLKINVX1 U21 ( .A(n123), .Y(n9) );
  CLKINVX1 U22 ( .A(n109), .Y(n12) );
  NAND2X1 U23 ( .A(n124), .B(n84), .Y(n113) );
  CLKINVX1 U24 ( .A(n137), .Y(n13) );
  NOR2X1 U25 ( .A(n13), .B(n84), .Y(n109) );
  CLKINVX1 U26 ( .A(n136), .Y(n20) );
  OAI22XL U27 ( .A0(n137), .A1(n17), .B0(n21), .B1(n12), .Y(n146) );
  OAI21X1 U28 ( .A0(n87), .A1(n8), .B0(n129), .Y(n141) );
  NAND2X1 U29 ( .A(n116), .B(n10), .Y(n129) );
  CLKINVX1 U30 ( .A(n93), .Y(n15) );
  OAI21XL U31 ( .A0(n119), .A1(n15), .B0(n118), .Y(n120) );
  OAI21XL U32 ( .A0(n125), .A1(n137), .B0(n124), .Y(n118) );
  NOR2X1 U34 ( .A(n10), .B(n85), .Y(n123) );
  CLKINVX1 U35 ( .A(n145), .Y(n85) );
  OAI22XL U36 ( .A0(n137), .A1(n113), .B0(n19), .B1(n9), .Y(n88) );
  CLKINVX1 U37 ( .A(n116), .Y(n83) );
  CLKINVX1 U38 ( .A(n131), .Y(n17) );
  CLKINVX1 U39 ( .A(n134), .Y(n14) );
  NOR2XL U40 ( .A(n125), .B(n87), .Y(n110) );
  CLKINVX1 U41 ( .A(n119), .Y(n11) );
  CLKINVX1 U42 ( .A(n103), .Y(n6) );
  OA21XL U43 ( .A0(n7), .A1(n15), .B0(n117), .Y(n102) );
  CLKINVX1 U45 ( .A(n105), .Y(n7) );
  OAI2BB1XL U46 ( .A0N(n103), .A1N(n124), .B0(n102), .Y(n104) );
  OAI22X1 U47 ( .A0(n10), .A1(n83), .B0(n4), .B1(n14), .Y(n112) );
  NOR4X1 U49 ( .A(n4), .B(addr[3]), .C(n21), .D(n86), .Y(n99) );
  XNOR2X1 U50 ( .A(addr[6]), .B(n5), .Y(n101) );
  AOI211X1 U53 ( .A0(n116), .A1(addr[6]), .B0(n115), .C0(n114), .Y(n128) );
  OAI222X1 U54 ( .A0(n111), .A1(n18), .B0(n110), .B1(n15), .C0(n20), .C1(n12), 
        .Y(n115) );
  OAI2BB2XL U55 ( .B0(n11), .B1(n113), .A0N(n21), .A1N(n112), .Y(n114) );
  OA21XL U56 ( .A0(n84), .A1(n3), .B0(n9), .Y(n111) );
  NAND2X1 U57 ( .A(n5), .B(n136), .Y(n133) );
  CLKINVX1 U59 ( .A(addr[6]), .Y(n19) );
  AOI211X1 U61 ( .A0(n131), .A1(n3), .B0(n92), .C0(n91), .Y(n95) );
  OAI221X1 U63 ( .A0(n21), .A1(n85), .B0(n18), .B1(n13), .C0(n102), .Y(n92) );
  OAI31X1 U64 ( .A0(n84), .A1(n87), .A2(n20), .B0(n90), .Y(n91) );
  AO21XL U66 ( .A0(n119), .A1(n129), .B0(addr[6]), .Y(n90) );
  NOR2X1 U67 ( .A(n87), .B(addr[3]), .Y(n145) );
  AOI21XL U68 ( .A0(addr[3]), .A1(n98), .B0(n97), .Y(n108) );
  OAI2BB1XL U69 ( .A0N(n86), .A1N(n124), .B0(n133), .Y(n98) );
  NAND3X1 U70 ( .A(n136), .B(n84), .C(n3), .Y(n117) );
  NOR2X1 U71 ( .A(addr[3]), .B(n3), .Y(n134) );
  OAI21X1 U72 ( .A0(n5), .A1(n142), .B0(n133), .Y(n138) );
  OAI22XL U73 ( .A0(n142), .A1(n83), .B0(n1), .B1(n132), .Y(n135) );
  AO21X1 U74 ( .A0(n139), .A1(n10), .B0(n138), .Y(n144) );
  OAI21XL U75 ( .A0(n2), .A1(n21), .B0(n15), .Y(n139) );
  OAI221X1 U76 ( .A0(n96), .A1(n86), .B0(n5), .B1(n95), .C0(n94), .Y(dout[1])
         );
  AOI2BB2X1 U77 ( .B0(n93), .B1(n112), .A0N(n133), .A1N(n6), .Y(n94) );
  OAI211X1 U78 ( .A0(n128), .A1(n86), .B0(n127), .C0(n126), .Y(dout[3]) );
  AOI32XL U79 ( .A0(n125), .A1(n1), .A2(n124), .B0(n123), .B1(n136), .Y(n126)
         );
  OAI31X1 U80 ( .A0(n122), .A1(n121), .A2(n120), .B0(n86), .Y(n127) );
  OAI221X1 U81 ( .A0(n3), .A1(n108), .B0(n107), .B1(n10), .C0(n106), .Y(
        dout[2]) );
  AOI32XL U82 ( .A0(n105), .A1(n86), .A2(n140), .B0(n2), .B1(n104), .Y(n106)
         );
  AOI211X1 U83 ( .A0(n101), .A1(n4), .B0(n100), .C0(n99), .Y(n107) );
  NAND2X1 U84 ( .A(n148), .B(n147), .Y(dout[4]) );
  AOI222XL U85 ( .A0(n136), .A1(n141), .B0(n3), .B1(n135), .C0(n134), .C1(n138), .Y(n148) );
  AOI222XL U86 ( .A0(n5), .A1(n146), .B0(n145), .B1(n144), .C0(n143), .C1(n86), 
        .Y(n147) );
  CLKINVX3 U87 ( .A(n3), .Y(n10) );
  CLKINVX3 U88 ( .A(addr[1]), .Y(n21) );
  CLKINVX3 U89 ( .A(addr[3]), .Y(n84) );
  CLKINVX3 U90 ( .A(n5), .Y(n86) );
  CLKINVX3 U91 ( .A(n4), .Y(n87) );
endmodule


module sbox8_11 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132;

  NAND2X2 U41 ( .A(addr[6]), .B(n6), .Y(n131) );
  NAND2X2 U48 ( .A(addr[4]), .B(n74), .Y(n123) );
  NAND2X2 U49 ( .A(n2), .B(n15), .Y(n87) );
  NAND2X2 U50 ( .A(addr[1]), .B(n16), .Y(n124) );
  NAND2X2 U54 ( .A(addr[2]), .B(n75), .Y(n116) );
  NAND2X2 U60 ( .A(addr[6]), .B(addr[1]), .Y(n105) );
  NAND2X2 U61 ( .A(n6), .B(n16), .Y(n108) );
  OAI32X1 U1 ( .A0(n16), .A1(addr[4]), .A2(n92), .B0(n115), .B1(n108), .Y(n96)
         );
  OAI31X1 U2 ( .A0(n123), .A1(addr[6]), .A2(n116), .B0(n109), .Y(n110) );
  OAI221X1 U3 ( .A0(n105), .A1(n87), .B0(addr[4]), .B1(n108), .C0(n86), .Y(n90) );
  NAND2X4 U4 ( .A(addr[4]), .B(n2), .Y(n115) );
  AOI222X1 U5 ( .A0(n88), .A1(addr[2]), .B0(n15), .B1(n10), .C0(n11), .C1(n92), 
        .Y(n114) );
  OAI222X1 U6 ( .A0(addr[2]), .A1(n126), .B0(n74), .B1(n125), .C0(n124), .C1(
        n123), .Y(n127) );
  AOI32XL U7 ( .A0(n9), .A1(n13), .A2(n2), .B0(n5), .B1(n117), .Y(n130) );
  OA21XL U8 ( .A0(n11), .A1(n75), .B0(n121), .Y(n78) );
  INVXL U9 ( .A(n119), .Y(n3) );
  INVX3 U10 ( .A(n2), .Y(n74) );
  BUFX4 U11 ( .A(addr[3]), .Y(n2) );
  CLKBUFX3 U12 ( .A(addr[5]), .Y(n1) );
  CLKINVX1 U13 ( .A(n108), .Y(n5) );
  CLKINVX1 U14 ( .A(n107), .Y(n12) );
  CLKINVX1 U15 ( .A(n93), .Y(n14) );
  NAND2X1 U16 ( .A(n74), .B(n15), .Y(n93) );
  NAND2X1 U17 ( .A(n11), .B(n75), .Y(n121) );
  OAI21XL U18 ( .A0(n115), .A1(n75), .B0(n107), .Y(n77) );
  OAI21X1 U19 ( .A0(n15), .A1(n75), .B0(n123), .Y(n88) );
  OAI31XL U20 ( .A0(n115), .A1(n6), .A2(n116), .B0(n118), .Y(n94) );
  CLKINVX1 U21 ( .A(n131), .Y(n4) );
  NAND2X1 U22 ( .A(n13), .B(n74), .Y(n107) );
  OAI22XL U23 ( .A0(n116), .A1(n123), .B0(n13), .B1(n115), .Y(n117) );
  OAI22XL U24 ( .A0(n123), .A1(n108), .B0(n131), .B1(n93), .Y(n95) );
  OAI2BB2XL U25 ( .B0(n115), .B1(n131), .A0N(n88), .A1N(n8), .Y(n89) );
  AOI211XL U26 ( .A0(n108), .A1(n105), .B0(n15), .C0(n121), .Y(n85) );
  CLKINVX1 U27 ( .A(n124), .Y(n9) );
  OAI22XL U28 ( .A0(n13), .A1(n123), .B0(n78), .B1(n87), .Y(n81) );
  NAND2BX2 U29 ( .AN(n78), .B(n74), .Y(n120) );
  NAND2XL U30 ( .A(n115), .B(n93), .Y(n104) );
  OAI2BB2XL U31 ( .B0(n106), .B1(n105), .A0N(n104), .A1N(n9), .Y(n111) );
  NOR2BXL U32 ( .AN(n123), .B(n103), .Y(n106) );
  NAND3X1 U33 ( .A(n104), .B(n6), .C(n13), .Y(n84) );
  AO21X1 U34 ( .A0(n13), .A1(n8), .B0(n101), .Y(n102) );
  OAI33X1 U35 ( .A0(n16), .A1(n74), .A2(n100), .B0(n11), .B1(n103), .B2(n124), 
        .Y(n101) );
  OA22XL U36 ( .A0(n107), .A1(n131), .B0(n120), .B1(n124), .Y(n98) );
  CLKINVX1 U37 ( .A(n125), .Y(n7) );
  OAI21XL U38 ( .A0(n9), .A1(n4), .B0(addr[4]), .Y(n86) );
  NAND2X1 U39 ( .A(n1), .B(n11), .Y(n100) );
  OAI221X1 U40 ( .A0(n124), .A1(n121), .B0(addr[1]), .B1(n120), .C0(n3), .Y(
        n128) );
  OAI31XL U42 ( .A0(n11), .A1(n6), .A2(n74), .B0(n118), .Y(n119) );
  NAND2X1 U43 ( .A(n8), .B(addr[2]), .Y(n125) );
  NAND4XL U44 ( .A(n4), .B(n1), .C(n2), .D(addr[2]), .Y(n109) );
  NAND3X1 U45 ( .A(n13), .B(n16), .C(n2), .Y(n118) );
  OAI21XL U46 ( .A0(n1), .A1(n87), .B0(n114), .Y(n76) );
  OAI22XL U47 ( .A0(n108), .A1(n120), .B0(n79), .B1(n100), .Y(n80) );
  AOI221XL U51 ( .A0(n4), .A1(n74), .B0(n8), .B1(n2), .C0(n91), .Y(n79) );
  NOR2X1 U52 ( .A(n1), .B(n2), .Y(n103) );
  NOR2X1 U53 ( .A(n87), .B(addr[6]), .Y(n91) );
  NOR2X1 U55 ( .A(n74), .B(n1), .Y(n92) );
  CLKINVX1 U56 ( .A(n100), .Y(n10) );
  OA21XL U57 ( .A0(n1), .A1(n115), .B0(n120), .Y(n132) );
  AOI221XL U58 ( .A0(n5), .A1(n2), .B0(n8), .B1(addr[4]), .C0(n122), .Y(n126)
         );
  OAI22XL U59 ( .A0(n2), .A1(n6), .B0(addr[4]), .B1(n131), .Y(n122) );
  OAI211X1 U62 ( .A0(addr[2]), .A1(n99), .B0(n98), .C0(n97), .Y(dout[2]) );
  AOI221XL U63 ( .A0(addr[2]), .A1(n96), .B0(n1), .B1(n95), .C0(n94), .Y(n97)
         );
  AOI221XL U64 ( .A0(n91), .A1(n1), .B0(n90), .B1(n75), .C0(n89), .Y(n99) );
  OAI211X1 U65 ( .A0(n132), .A1(n131), .B0(n130), .C0(n129), .Y(dout[4]) );
  AOI222XL U66 ( .A0(n128), .A1(n15), .B0(n1), .B1(n127), .C0(n12), .C1(n8), 
        .Y(n129) );
  OAI211X1 U67 ( .A0(addr[1]), .A1(n114), .B0(n113), .C0(n112), .Y(dout[3]) );
  AOI221XL U68 ( .A0(n111), .A1(n11), .B0(n12), .B1(n5), .C0(n110), .Y(n112)
         );
  AOI2BB2XL U69 ( .B0(n102), .B1(n15), .A0N(n115), .A1N(n125), .Y(n113) );
  NAND4BX1 U70 ( .AN(n85), .B(n84), .C(n83), .D(n82), .Y(dout[1]) );
  AOI221XL U71 ( .A0(n4), .A1(n81), .B0(n14), .B1(n7), .C0(n80), .Y(n82) );
  AOI22X1 U72 ( .A0(n8), .A1(n77), .B0(n9), .B1(n76), .Y(n83) );
  CLKINVX3 U73 ( .A(addr[1]), .Y(n6) );
  CLKINVX3 U74 ( .A(n105), .Y(n8) );
  CLKINVX3 U75 ( .A(addr[2]), .Y(n11) );
  CLKINVX3 U76 ( .A(n116), .Y(n13) );
  CLKINVX3 U77 ( .A(addr[4]), .Y(n15) );
  CLKINVX3 U78 ( .A(addr[6]), .Y(n16) );
  CLKINVX3 U79 ( .A(n1), .Y(n75) );
endmodule


module crp_11 ( P, R, K_sub );
  output [1:32] P;
  input [1:32] R;
  input [1:48] K_sub;
  wire   n1;
  wire   [1:48] X;

  sbox1_11 u0 ( .addr(X[1:6]), .dout({P[9], P[17], P[23], P[31]}) );
  sbox2_11 u1 ( .addr({X[7], n1, X[9:12]}), .dout({P[13], P[28], P[2], P[18]})
         );
  sbox3_11 u2 ( .addr(X[13:18]), .dout({P[24], P[16], P[30], P[6]}) );
  sbox4_11 u3 ( .addr(X[19:24]), .dout({P[26], P[20], P[10], P[1]}) );
  sbox5_11 u4 ( .addr(X[25:30]), .dout({P[8], P[14], P[25], P[3]}) );
  sbox6_11 u5 ( .addr(X[31:36]), .dout({P[4], P[29], P[11], P[19]}) );
  sbox7_11 u6 ( .addr(X[37:42]), .dout({P[32], P[12], P[22], P[7]}) );
  sbox8_11 u7 ( .addr(X[43:48]), .dout({P[5], P[27], P[15], P[21]}) );
  XOR2X1 U1 ( .A(R[1]), .B(K_sub[2]), .Y(X[2]) );
  CLKXOR2X4 U2 ( .A(R[29]), .B(K_sub[42]), .Y(X[42]) );
  CLKXOR2X4 U3 ( .A(R[5]), .B(K_sub[6]), .Y(X[6]) );
  CLKXOR2X4 U4 ( .A(R[16]), .B(K_sub[25]), .Y(X[25]) );
  CLKXOR2X4 U5 ( .A(R[8]), .B(K_sub[11]), .Y(X[11]) );
  CLKXOR2X4 U6 ( .A(R[22]), .B(K_sub[33]), .Y(X[33]) );
  CLKXOR2X4 U7 ( .A(R[16]), .B(K_sub[23]), .Y(X[23]) );
  CLKXOR2X4 U8 ( .A(R[10]), .B(K_sub[15]), .Y(X[15]) );
  XNOR2X1 U9 ( .A(R[5]), .B(K_sub[8]), .Y(X[8]) );
  INVX3 U10 ( .A(X[8]), .Y(n1) );
  CLKXOR2X4 U11 ( .A(R[20]), .B(K_sub[31]), .Y(X[31]) );
  CLKXOR2X4 U12 ( .A(R[31]), .B(K_sub[46]), .Y(X[46]) );
  CLKXOR2X4 U13 ( .A(R[29]), .B(K_sub[44]), .Y(X[44]) );
  CLKXOR2X4 U14 ( .A(R[12]), .B(K_sub[19]), .Y(X[19]) );
  CLKXOR2X4 U15 ( .A(R[26]), .B(K_sub[39]), .Y(X[39]) );
  CLKXOR2X4 U16 ( .A(R[20]), .B(K_sub[29]), .Y(X[29]) );
  CLKXOR2X2 U17 ( .A(R[4]), .B(K_sub[5]), .Y(X[5]) );
  CLKXOR2X2 U18 ( .A(R[15]), .B(K_sub[22]), .Y(X[22]) );
  CLKXOR2X2 U19 ( .A(R[24]), .B(K_sub[35]), .Y(X[35]) );
  CLKXOR2X2 U20 ( .A(R[21]), .B(K_sub[30]), .Y(X[30]) );
  CLKXOR2X2 U21 ( .A(R[12]), .B(K_sub[17]), .Y(X[17]) );
  CLKXOR2X2 U22 ( .A(R[32]), .B(K_sub[1]), .Y(X[1]) );
  CLKXOR2X2 U23 ( .A(R[13]), .B(K_sub[20]), .Y(X[20]) );
  CLKXOR2X2 U24 ( .A(R[18]), .B(K_sub[27]), .Y(X[27]) );
  CLKXOR2X2 U25 ( .A(R[8]), .B(K_sub[13]), .Y(X[13]) );
  CLKXOR2X2 U26 ( .A(R[4]), .B(K_sub[7]), .Y(X[7]) );
  CLKXOR2X2 U27 ( .A(R[24]), .B(K_sub[37]), .Y(X[37]) );
  CLKXOR2X2 U28 ( .A(R[28]), .B(K_sub[43]), .Y(X[43]) );
  CLKXOR2X2 U29 ( .A(R[1]), .B(K_sub[48]), .Y(X[48]) );
  CLKXOR2X2 U30 ( .A(R[17]), .B(K_sub[24]), .Y(X[24]) );
  CLKXOR2X2 U31 ( .A(R[9]), .B(K_sub[12]), .Y(X[12]) );
  CLKXOR2X2 U32 ( .A(R[13]), .B(K_sub[18]), .Y(X[18]) );
  CLKXOR2X2 U33 ( .A(R[25]), .B(K_sub[36]), .Y(X[36]) );
  XOR2X1 U34 ( .A(R[23]), .B(K_sub[34]), .Y(X[34]) );
  XOR2X1 U35 ( .A(R[9]), .B(K_sub[14]), .Y(X[14]) );
  XOR2X1 U36 ( .A(R[30]), .B(K_sub[45]), .Y(X[45]) );
  XOR2X1 U37 ( .A(R[21]), .B(K_sub[32]), .Y(X[32]) );
  XOR2X1 U38 ( .A(R[25]), .B(K_sub[38]), .Y(X[38]) );
  XOR2X1 U39 ( .A(R[27]), .B(K_sub[40]), .Y(X[40]) );
  XOR2X1 U40 ( .A(R[3]), .B(K_sub[4]), .Y(X[4]) );
  XOR2X1 U41 ( .A(R[11]), .B(K_sub[16]), .Y(X[16]) );
  XOR2X1 U42 ( .A(R[7]), .B(K_sub[10]), .Y(X[10]) );
  XOR2X1 U43 ( .A(R[14]), .B(K_sub[21]), .Y(X[21]) );
  XOR2X1 U44 ( .A(R[6]), .B(K_sub[9]), .Y(X[9]) );
  XOR2X1 U45 ( .A(R[2]), .B(K_sub[3]), .Y(X[3]) );
  XOR2X1 U46 ( .A(R[28]), .B(K_sub[41]), .Y(X[41]) );
  XOR2X1 U47 ( .A(R[17]), .B(K_sub[26]), .Y(X[26]) );
  XOR2X1 U48 ( .A(R[32]), .B(K_sub[47]), .Y(X[47]) );
  XOR2X1 U49 ( .A(R[19]), .B(K_sub[28]), .Y(X[28]) );
endmodule


module sbox1_10 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127;

  OAI222X4 U13 ( .A0(addr[5]), .A1(n101), .B0(n1), .B1(n100), .C0(n99), .C1(
        n10), .Y(dout[3]) );
  OAI21X2 U42 ( .A0(n4), .A1(n112), .B0(n106), .Y(n123) );
  NAND2X2 U44 ( .A(addr[6]), .B(n72), .Y(n115) );
  NAND2X2 U48 ( .A(addr[1]), .B(n13), .Y(n114) );
  OAI22X2 U49 ( .A0(n6), .A1(n71), .B0(addr[5]), .B1(n120), .Y(n85) );
  NAND2X2 U50 ( .A(n3), .B(n6), .Y(n120) );
  NOR2X2 U51 ( .A(n6), .B(n3), .Y(n124) );
  NOR2X2 U56 ( .A(n109), .B(n3), .Y(n93) );
  NAND2X2 U57 ( .A(addr[1]), .B(addr[6]), .Y(n109) );
  NAND2X2 U59 ( .A(n72), .B(n13), .Y(n112) );
  NOR2X1 U1 ( .A(n114), .B(n120), .Y(n104) );
  AOI221X4 U2 ( .A0(n12), .A1(n90), .B0(n4), .B1(n93), .C0(n102), .Y(n79) );
  NOR3X1 U3 ( .A(n2), .B(addr[6]), .C(n10), .Y(n102) );
  BUFX4 U4 ( .A(addr[4]), .Y(n2) );
  CLKBUFX3 U5 ( .A(addr[2]), .Y(n1) );
  OAI32X1 U6 ( .A0(n112), .A1(n2), .A2(n4), .B0(n115), .B1(n113), .Y(n80) );
  NOR2BXL U7 ( .AN(n118), .B(n1), .Y(n122) );
  CLKBUFX3 U8 ( .A(addr[2]), .Y(n4) );
  OAI221X4 U9 ( .A0(addr[5]), .A1(n127), .B0(n126), .B1(n71), .C0(n125), .Y(
        dout[4]) );
  OAI221X4 U10 ( .A0(n88), .A1(n71), .B0(addr[5]), .B1(n87), .C0(n86), .Y(
        dout[2]) );
  OA21XL U11 ( .A0(n95), .A1(n115), .B0(n107), .Y(n119) );
  AOI222XL U12 ( .A0(n12), .A1(n1), .B0(n2), .B1(n110), .C0(n69), .C1(n10), 
        .Y(n111) );
  AOI2BB2X1 U14 ( .B0(n2), .B1(n69), .A0N(addr[4]), .A1N(n115), .Y(n91) );
  BUFX4 U15 ( .A(addr[3]), .Y(n3) );
  CLKINVX1 U16 ( .A(n112), .Y(n12) );
  CLKINVX1 U17 ( .A(n113), .Y(n7) );
  NAND2BX1 U18 ( .AN(n104), .B(n119), .Y(n84) );
  CLKXOR2X2 U19 ( .A(n8), .B(n10), .Y(n90) );
  NOR2X1 U20 ( .A(n6), .B(n8), .Y(n118) );
  OAI21XL U21 ( .A0(n8), .A1(n114), .B0(n91), .Y(n92) );
  NAND2X1 U22 ( .A(n93), .B(n6), .Y(n107) );
  NAND2X1 U23 ( .A(n10), .B(n8), .Y(n113) );
  OAI211X1 U24 ( .A0(n6), .A1(n114), .B0(n108), .C0(n107), .Y(n89) );
  CLKINVX1 U25 ( .A(n109), .Y(n69) );
  NAND2X1 U26 ( .A(n124), .B(n70), .Y(n108) );
  CLKINVX1 U27 ( .A(n114), .Y(n11) );
  CLKINVX1 U28 ( .A(n115), .Y(n70) );
  CLKINVX1 U29 ( .A(n95), .Y(n9) );
  AO22X1 U30 ( .A0(n90), .A1(n70), .B0(n8), .B1(n123), .Y(n76) );
  OAI31X1 U31 ( .A0(n10), .A1(n3), .A2(n72), .B0(n103), .Y(n105) );
  AOI31XL U32 ( .A0(n72), .A1(n10), .A2(n2), .B0(n102), .Y(n103) );
  CLKINVX1 U33 ( .A(addr[6]), .Y(n13) );
  AOI211X1 U34 ( .A0(n5), .A1(n4), .B0(n117), .C0(n116), .Y(n126) );
  CLKINVX1 U35 ( .A(n108), .Y(n5) );
  AOI211X1 U36 ( .A0(n115), .A1(n114), .B0(n113), .C0(n2), .Y(n116) );
  OAI22X1 U37 ( .A0(n120), .A1(n112), .B0(n111), .B1(n8), .Y(n117) );
  AOI211X1 U38 ( .A0(n69), .A1(n118), .B0(n81), .C0(n80), .Y(n88) );
  OAI22X1 U39 ( .A0(n91), .A1(n10), .B0(n3), .B1(n106), .Y(n81) );
  CLKINVX3 U40 ( .A(addr[5]), .Y(n71) );
  NAND2X1 U41 ( .A(n3), .B(n71), .Y(n95) );
  NAND2X1 U43 ( .A(n11), .B(n1), .Y(n106) );
  XOR2X1 U45 ( .A(n82), .B(n2), .Y(n83) );
  NAND2X1 U46 ( .A(n1), .B(n3), .Y(n82) );
  OAI22XL U47 ( .A0(n3), .A1(n72), .B0(n8), .B1(n112), .Y(n94) );
  AOI211XL U52 ( .A0(n98), .A1(n8), .B0(n97), .C0(n104), .Y(n99) );
  OAI22XL U53 ( .A0(n96), .A1(n6), .B0(n95), .B1(n109), .Y(n97) );
  OAI22XL U54 ( .A0(n13), .A1(n71), .B0(n2), .B1(addr[1]), .Y(n98) );
  AOI221XL U55 ( .A0(n9), .A1(addr[6]), .B0(addr[5]), .B1(n94), .C0(n93), .Y(
        n96) );
  OAI21XL U58 ( .A0(addr[1]), .A1(n120), .B0(n119), .Y(n121) );
  AOI221XL U60 ( .A0(n12), .A1(n118), .B0(n93), .B1(n71), .C0(n75), .Y(n78) );
  OAI31X1 U61 ( .A0(n71), .A1(n2), .A2(n74), .B0(n73), .Y(n75) );
  OA21XL U62 ( .A0(n3), .A1(n13), .B0(n109), .Y(n74) );
  OAI21XL U63 ( .A0(n124), .A1(n85), .B0(n11), .Y(n73) );
  OAI21XL U64 ( .A0(n1), .A1(n72), .B0(n109), .Y(n110) );
  INVX4 U65 ( .A(n4), .Y(n10) );
  AOI222XL U66 ( .A0(n124), .A1(n123), .B0(n122), .B1(addr[6]), .C0(n1), .C1(
        n121), .Y(n125) );
  NOR4BBX1 U67 ( .AN(n107), .BN(n106), .C(n105), .D(n104), .Y(n127) );
  AOI222XL U68 ( .A0(n12), .A1(n90), .B0(n89), .B1(n10), .C0(n123), .C1(n6), 
        .Y(n101) );
  AOI2BB2XL U69 ( .B0(addr[5]), .B1(n92), .A0N(n120), .A1N(addr[1]), .Y(n100)
         );
  AOI32X1 U70 ( .A0(n4), .A1(n85), .A2(n12), .B0(n84), .B1(n10), .Y(n86) );
  AOI222XL U71 ( .A0(n124), .A1(n72), .B0(n83), .B1(addr[1]), .C0(n7), .C1(n13), .Y(n87) );
  OAI221X1 U72 ( .A0(n79), .A1(n71), .B0(n4), .B1(n78), .C0(n77), .Y(dout[1])
         );
  AOI32XL U73 ( .A0(addr[6]), .A1(n85), .A2(n1), .B0(n76), .B1(n71), .Y(n77)
         );
  CLKINVX3 U74 ( .A(n2), .Y(n6) );
  CLKINVX3 U75 ( .A(n3), .Y(n8) );
  CLKINVX3 U76 ( .A(addr[1]), .Y(n72) );
endmodule


module sbox2_10 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147;

  NAND2X2 U55 ( .A(n2), .B(n81), .Y(n136) );
  NAND2X2 U57 ( .A(addr[2]), .B(n15), .Y(n104) );
  NAND2X2 U60 ( .A(addr[5]), .B(addr[2]), .Y(n132) );
  NOR2X2 U61 ( .A(n7), .B(n4), .Y(n101) );
  NAND2X2 U62 ( .A(n6), .B(n13), .Y(n146) );
  NAND2X2 U63 ( .A(n3), .B(n83), .Y(n124) );
  NAND2X2 U64 ( .A(addr[6]), .B(n6), .Y(n122) );
  NAND2X2 U67 ( .A(n3), .B(n2), .Y(n133) );
  AOI222XL U1 ( .A0(n9), .A1(n8), .B0(n88), .B1(n83), .C0(n140), .C1(n4), .Y(
        n89) );
  CLKINVX1 U2 ( .A(n121), .Y(n7) );
  OAI211X4 U3 ( .A0(n147), .A1(n146), .B0(n145), .C0(n144), .Y(dout[4]) );
  CLKINVX1 U4 ( .A(addr[5]), .Y(n1) );
  INVX3 U5 ( .A(addr[5]), .Y(n15) );
  NAND3XL U6 ( .A(n98), .B(n97), .C(n96), .Y(dout[1]) );
  NAND2X1 U7 ( .A(addr[1]), .B(addr[6]), .Y(n121) );
  CLKINVX2 U8 ( .A(addr[1]), .Y(n6) );
  OAI221X1 U9 ( .A0(addr[1]), .A1(n136), .B0(n133), .B1(n6), .C0(n87), .Y(n95)
         );
  NOR2X1 U10 ( .A(n104), .B(n2), .Y(n141) );
  NOR2X1 U11 ( .A(n124), .B(n2), .Y(n140) );
  CLKBUFX4 U12 ( .A(addr[4]), .Y(n2) );
  NAND2X4 U13 ( .A(addr[1]), .B(n13), .Y(n114) );
  INVX3 U14 ( .A(addr[6]), .Y(n13) );
  NAND2XL U15 ( .A(n102), .B(n81), .Y(n109) );
  AOI211XL U16 ( .A0(n16), .A1(n95), .B0(n94), .C0(n93), .Y(n96) );
  AOI2BB2X1 U17 ( .B0(n15), .B1(n82), .A0N(n104), .A1N(n136), .Y(n117) );
  NOR3BXL U18 ( .AN(n135), .B(n134), .C(n9), .Y(n147) );
  BUFX4 U19 ( .A(addr[3]), .Y(n3) );
  NAND2X1 U20 ( .A(n9), .B(n7), .Y(n113) );
  CLKINVX1 U21 ( .A(n146), .Y(n4) );
  CLKINVX1 U22 ( .A(n115), .Y(n9) );
  CLKINVX1 U23 ( .A(n122), .Y(n5) );
  OAI31X1 U24 ( .A0(n124), .A1(n13), .A2(n15), .B0(n123), .Y(n128) );
  OAI21XL U25 ( .A0(n15), .A1(n6), .B0(n140), .Y(n123) );
  OAI22X1 U26 ( .A0(n122), .A1(n124), .B0(n101), .B1(n132), .Y(n84) );
  INVX1 U27 ( .A(n114), .Y(n8) );
  OAI22X1 U28 ( .A0(n122), .A1(n81), .B0(n10), .B1(n121), .Y(n129) );
  NAND3X1 U29 ( .A(n10), .B(n15), .C(n6), .Y(n111) );
  NAND2X1 U30 ( .A(n81), .B(n10), .Y(n115) );
  OAI21XL U31 ( .A0(n83), .A1(n133), .B0(n135), .Y(n85) );
  OAI22XL U32 ( .A0(n117), .A1(n146), .B0(n116), .B1(n132), .Y(n118) );
  AOI222XL U33 ( .A0(n8), .A1(n115), .B0(n11), .B1(n13), .C0(n9), .C1(n4), .Y(
        n116) );
  CLKINVX1 U34 ( .A(n104), .Y(n14) );
  OAI2BB2XL U35 ( .B0(n114), .B1(n135), .A0N(n126), .A1N(n11), .Y(n106) );
  OAI21XL U36 ( .A0(n112), .A1(n114), .B0(n111), .Y(n120) );
  OAI21XL U37 ( .A0(n133), .A1(n114), .B0(n113), .Y(n119) );
  CLKINVX1 U38 ( .A(n124), .Y(n82) );
  CLKINVX1 U39 ( .A(n136), .Y(n12) );
  CLKINVX1 U40 ( .A(n133), .Y(n11) );
  CLKINVX1 U41 ( .A(n132), .Y(n16) );
  AOI2BB1X1 U42 ( .A0N(n126), .A1N(n125), .B0(n136), .Y(n127) );
  OAI22XL U43 ( .A0(n104), .A1(n114), .B0(n101), .B1(n132), .Y(n102) );
  AO21XL U44 ( .A0(n83), .A1(n12), .B0(n141), .Y(n86) );
  AO21X1 U45 ( .A0(n81), .A1(n14), .B0(n140), .Y(n142) );
  NAND3X1 U46 ( .A(n83), .B(n10), .C(addr[5]), .Y(n135) );
  OAI22X1 U47 ( .A0(addr[5]), .A1(n121), .B0(n122), .B1(n15), .Y(n126) );
  AOI2BB1X1 U48 ( .A0N(n3), .A1N(n1), .B0(n12), .Y(n112) );
  NOR3X1 U49 ( .A(addr[1]), .B(addr[2]), .C(n15), .Y(n125) );
  AOI2BB1XL U50 ( .A0N(n92), .A1N(n91), .B0(addr[5]), .Y(n93) );
  OAI22XL U51 ( .A0(n117), .A1(n114), .B0(n89), .B1(n1), .Y(n94) );
  OAI31XL U52 ( .A0(n114), .A1(n2), .A2(n81), .B0(n90), .Y(n91) );
  OAI21XL U53 ( .A0(n11), .A1(n82), .B0(n5), .Y(n90) );
  NAND2X1 U54 ( .A(n8), .B(n2), .Y(n137) );
  OAI31XL U56 ( .A0(n101), .A1(n3), .A2(addr[2]), .B0(n113), .Y(n92) );
  OAI211X1 U58 ( .A0(n139), .A1(n15), .B0(n138), .C0(n137), .Y(n143) );
  NAND3X1 U59 ( .A(n10), .B(n15), .C(addr[6]), .Y(n138) );
  AOI2BB2X1 U65 ( .B0(n5), .B1(n81), .A0N(n6), .A1N(n136), .Y(n139) );
  OAI22XL U66 ( .A0(addr[5]), .A1(n133), .B0(n3), .B1(n132), .Y(n134) );
  OAI2BB2XL U68 ( .B0(n112), .B1(n122), .A0N(n1), .A1N(n99), .Y(n100) );
  OAI211X1 U69 ( .A0(n146), .A1(n2), .B0(n137), .C0(n113), .Y(n99) );
  NAND3X1 U70 ( .A(n5), .B(n10), .C(n3), .Y(n87) );
  AOI2BB2XL U71 ( .B0(n3), .B1(n105), .A0N(n137), .A1N(n132), .Y(n108) );
  OAI211XL U72 ( .A0(n104), .A1(n146), .B0(n103), .C0(n111), .Y(n105) );
  NAND3XL U73 ( .A(addr[5]), .B(n10), .C(n7), .Y(n103) );
  OAI22XL U74 ( .A0(n3), .A1(n114), .B0(n13), .B1(n115), .Y(n88) );
  NAND4X1 U75 ( .A(n110), .B(n109), .C(n108), .D(n107), .Y(dout[2]) );
  AOI32XL U76 ( .A0(addr[1]), .A1(addr[2]), .A2(n12), .B0(n100), .B1(n83), .Y(
        n110) );
  AOI221XL U77 ( .A0(n125), .A1(addr[4]), .B0(n141), .B1(n5), .C0(n106), .Y(
        n107) );
  AOI33XL U78 ( .A0(n5), .A1(n14), .A2(n2), .B0(n16), .B1(n146), .B2(n3), .Y(
        n145) );
  AOI222XL U79 ( .A0(n143), .A1(n83), .B0(n7), .B1(n142), .C0(n8), .C1(n141), 
        .Y(n144) );
  AOI32XL U80 ( .A0(n14), .A1(n6), .A2(n9), .B0(n4), .B1(n86), .Y(n97) );
  AOI22X1 U81 ( .A0(n7), .A1(n85), .B0(n2), .B1(n84), .Y(n98) );
  NAND2X1 U82 ( .A(n131), .B(n130), .Y(dout[3]) );
  AOI221XL U83 ( .A0(n120), .A1(n83), .B0(addr[2]), .B1(n119), .C0(n118), .Y(
        n131) );
  AOI211X1 U84 ( .A0(n14), .A1(n129), .B0(n128), .C0(n127), .Y(n130) );
  CLKINVX3 U85 ( .A(n2), .Y(n10) );
  CLKINVX3 U86 ( .A(n3), .Y(n81) );
  CLKINVX3 U87 ( .A(addr[2]), .Y(n83) );
endmodule


module sbox3_10 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134;

  NOR2X2 U35 ( .A(n14), .B(addr[3]), .Y(n109) );
  NOR2X2 U50 ( .A(addr[1]), .B(addr[6]), .Y(n108) );
  NOR2X2 U52 ( .A(n16), .B(n3), .Y(n88) );
  NOR2X2 U56 ( .A(n16), .B(n8), .Y(n95) );
  NOR2X1 U1 ( .A(n14), .B(n16), .Y(n107) );
  OAI221X1 U2 ( .A0(n125), .A1(n14), .B0(n4), .B1(addr[1]), .C0(n77), .Y(n105)
         );
  INVXL U3 ( .A(n2), .Y(n1) );
  NOR2X1 U4 ( .A(n76), .B(n4), .Y(n92) );
  NOR2X1 U5 ( .A(n15), .B(n4), .Y(n122) );
  NOR2X1 U6 ( .A(n77), .B(n4), .Y(n96) );
  CLKBUFX3 U7 ( .A(addr[2]), .Y(n4) );
  INVX1 U8 ( .A(addr[2]), .Y(n2) );
  NOR2X1 U9 ( .A(n4), .B(n3), .Y(n111) );
  BUFX4 U10 ( .A(addr[4]), .Y(n3) );
  OAI33X1 U11 ( .A0(n15), .A1(n126), .A2(n8), .B0(n14), .B1(n95), .B2(n120), 
        .Y(n80) );
  INVX3 U12 ( .A(n4), .Y(n8) );
  OAI221X1 U13 ( .A0(addr[5]), .A1(n91), .B0(n90), .B1(n78), .C0(n89), .Y(
        dout[1]) );
  NOR2X4 U14 ( .A(n79), .B(n20), .Y(n125) );
  NOR2X4 U15 ( .A(addr[3]), .B(n3), .Y(n131) );
  NOR2X4 U16 ( .A(n20), .B(addr[6]), .Y(n126) );
  INVX3 U17 ( .A(addr[1]), .Y(n20) );
  NAND2XL U18 ( .A(n95), .B(n125), .Y(n133) );
  OAI211XL U19 ( .A0(n3), .A1(n9), .B0(n129), .C0(n128), .Y(n130) );
  NAND4XL U20 ( .A(n115), .B(n114), .C(n113), .D(n112), .Y(n116) );
  CLKINVX1 U21 ( .A(n133), .Y(n7) );
  INVX1 U22 ( .A(n125), .Y(n17) );
  CLKINVX1 U23 ( .A(n107), .Y(n12) );
  NAND2X1 U24 ( .A(n76), .B(n13), .Y(n123) );
  CLKINVX1 U25 ( .A(n87), .Y(n13) );
  CLKINVX1 U26 ( .A(n121), .Y(n5) );
  CLKINVX1 U27 ( .A(n120), .Y(n18) );
  CLKINVX1 U28 ( .A(n115), .Y(n6) );
  CLKINVX1 U29 ( .A(n108), .Y(n77) );
  NOR2X1 U30 ( .A(n76), .B(n8), .Y(n104) );
  NOR2X1 U31 ( .A(n17), .B(n8), .Y(n110) );
  INVX1 U32 ( .A(n126), .Y(n19) );
  AOI21X1 U33 ( .A0(n16), .A1(n8), .B0(n95), .Y(n121) );
  OAI21XL U34 ( .A0(n111), .A1(n131), .B0(n125), .Y(n83) );
  CLKINVX1 U36 ( .A(n82), .Y(n76) );
  NOR2X1 U37 ( .A(n19), .B(n14), .Y(n87) );
  NOR2X1 U38 ( .A(n125), .B(n108), .Y(n120) );
  OAI21XL U39 ( .A0(n110), .A1(n92), .B0(n131), .Y(n101) );
  NAND2X1 U40 ( .A(n104), .B(n88), .Y(n115) );
  CLKINVX1 U41 ( .A(n88), .Y(n15) );
  CLKINVX1 U42 ( .A(n92), .Y(n9) );
  CLKINVX1 U43 ( .A(n111), .Y(n10) );
  CLKINVX1 U44 ( .A(n122), .Y(n11) );
  OR2X1 U45 ( .A(n104), .B(n96), .Y(n127) );
  OAI221X1 U46 ( .A0(n19), .A1(n10), .B0(n8), .B1(n13), .C0(n94), .Y(n99) );
  AOI221XL U47 ( .A0(n96), .A1(n3), .B0(n93), .B1(n14), .C0(n7), .Y(n94) );
  OAI21XL U48 ( .A0(n8), .A1(n77), .B0(n9), .Y(n93) );
  XNOR2X1 U49 ( .A(addr[5]), .B(addr[3]), .Y(n103) );
  CLKINVX1 U51 ( .A(addr[5]), .Y(n78) );
  OAI221X1 U53 ( .A0(n77), .A1(n10), .B0(n17), .B1(n15), .C0(n106), .Y(n117)
         );
  AOI221XL U54 ( .A0(addr[3]), .A1(n105), .B0(n104), .B1(n131), .C0(n7), .Y(
        n106) );
  CLKINVX1 U55 ( .A(addr[6]), .Y(n79) );
  NAND3X1 U57 ( .A(n4), .B(n20), .C(n109), .Y(n114) );
  NOR2X1 U58 ( .A(n79), .B(addr[1]), .Y(n82) );
  AOI32XL U59 ( .A0(n8), .A1(n16), .A2(n125), .B0(n124), .B1(n79), .Y(n129) );
  AOI22XL U60 ( .A0(n3), .A1(n127), .B0(n126), .B1(n131), .Y(n128) );
  OAI22XL U61 ( .A0(n3), .A1(n2), .B0(n4), .B1(n12), .Y(n124) );
  AOI222XL U62 ( .A0(n111), .A1(n126), .B0(n110), .B1(n16), .C0(n109), .C1(
        n108), .Y(n112) );
  OAI211XL U63 ( .A0(n107), .A1(n131), .B0(n2), .C0(addr[6]), .Y(n113) );
  OAI21XL U64 ( .A0(n1), .A1(addr[1]), .B0(n19), .Y(n81) );
  AOI221XL U65 ( .A0(n87), .A1(n16), .B0(n88), .B1(n126), .C0(n86), .Y(n90) );
  OAI211X1 U66 ( .A0(n85), .A1(n8), .B0(n84), .C0(n83), .Y(n86) );
  AOI222XL U67 ( .A0(n82), .A1(n16), .B0(n108), .B1(n107), .C0(n131), .C1(n20), 
        .Y(n85) );
  OAI21XL U68 ( .A0(n92), .A1(n7), .B0(addr[4]), .Y(n84) );
  AOI221XL U69 ( .A0(n126), .A1(n5), .B0(addr[3]), .B1(n127), .C0(n97), .Y(n98) );
  OAI22X1 U70 ( .A0(n17), .A1(n11), .B0(n12), .B1(n76), .Y(n97) );
  OAI211X1 U71 ( .A0(n77), .A1(n11), .B0(n119), .C0(n118), .Y(dout[3]) );
  AOI32XL U72 ( .A0(n126), .A1(n4), .A2(n103), .B0(n109), .B1(n110), .Y(n119)
         );
  AOI22XL U73 ( .A0(n117), .A1(n78), .B0(addr[5]), .B1(n116), .Y(n118) );
  AOI221XL U74 ( .A0(n122), .A1(n126), .B0(n96), .B1(n109), .C0(n6), .Y(n89)
         );
  AOI221XL U75 ( .A0(n131), .A1(n81), .B0(n95), .B1(n123), .C0(n80), .Y(n91)
         );
  NAND4X1 U76 ( .A(n102), .B(n114), .C(n101), .D(n100), .Y(dout[2]) );
  NAND3XL U77 ( .A(n3), .B(n125), .C(n103), .Y(n102) );
  AOI2BB2XL U78 ( .B0(addr[5]), .B1(n99), .A0N(addr[5]), .A1N(n98), .Y(n100)
         );
  OAI221X1 U79 ( .A0(n134), .A1(n78), .B0(n3), .B1(n133), .C0(n132), .Y(
        dout[4]) );
  AOI32XL U80 ( .A0(n131), .A1(n79), .A2(n1), .B0(n130), .B1(n78), .Y(n132) );
  AOI222XL U81 ( .A0(n5), .A1(n123), .B0(n122), .B1(addr[1]), .C0(n121), .C1(
        n18), .Y(n134) );
  CLKINVX3 U82 ( .A(n3), .Y(n14) );
  CLKINVX3 U83 ( .A(addr[3]), .Y(n16) );
endmodule


module sbox4_10 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126;

  OAI32X4 U12 ( .A0(n16), .A1(n2), .A2(addr[2]), .B0(n72), .B1(n108), .Y(n123)
         );
  OAI222X4 U20 ( .A0(addr[2]), .A1(n92), .B0(n106), .B1(n91), .C0(n90), .C1(n9), .Y(dout[2]) );
  OAI222X4 U33 ( .A0(addr[4]), .A1(n106), .B0(n15), .B1(n108), .C0(n2), .C1(
        n118), .Y(n83) );
  NAND2X2 U34 ( .A(addr[4]), .B(n2), .Y(n108) );
  NOR2X2 U43 ( .A(n6), .B(addr[4]), .Y(n113) );
  NOR2X2 U45 ( .A(n72), .B(n2), .Y(n111) );
  NAND2X2 U51 ( .A(n15), .B(n12), .Y(n118) );
  NOR2X2 U52 ( .A(n71), .B(addr[5]), .Y(n97) );
  NAND2X2 U53 ( .A(addr[6]), .B(addr[1]), .Y(n85) );
  NAND2X2 U54 ( .A(addr[1]), .B(n12), .Y(n116) );
  NOR2X2 U55 ( .A(n115), .B(n72), .Y(n121) );
  NAND2X2 U56 ( .A(n6), .B(n71), .Y(n115) );
  NAND2X2 U57 ( .A(addr[5]), .B(n71), .Y(n96) );
  NAND2X2 U58 ( .A(addr[6]), .B(n15), .Y(n106) );
  OAI222X1 U1 ( .A0(n16), .A1(n85), .B0(n97), .B1(n116), .C0(n71), .C1(n118), 
        .Y(n73) );
  CLKINVX1 U2 ( .A(n116), .Y(n11) );
  OAI31X4 U3 ( .A0(n118), .A1(n72), .A2(n71), .B0(n117), .Y(n119) );
  CLKINVX1 U4 ( .A(n6), .Y(n1) );
  CLKBUFX3 U5 ( .A(addr[3]), .Y(n2) );
  OAI221X1 U6 ( .A0(addr[2]), .A1(n80), .B0(n118), .B1(n105), .C0(n79), .Y(
        dout[1]) );
  INVX4 U7 ( .A(addr[5]), .Y(n72) );
  OAI31X1 U8 ( .A0(n108), .A1(addr[5]), .A2(n13), .B0(n107), .Y(n109) );
  AOI222XL U9 ( .A0(n71), .A1(n12), .B0(n113), .B1(n15), .C0(addr[1]), .C1(n6), 
        .Y(n114) );
  OAI222X1 U10 ( .A0(addr[1]), .A1(n84), .B0(n85), .B1(n74), .C0(n6), .C1(n107), .Y(n75) );
  NAND2XL U11 ( .A(n1), .B(addr[5]), .Y(n84) );
  AOI211XL U13 ( .A0(n83), .A1(n72), .B0(n82), .C0(n5), .Y(n92) );
  NAND2XL U14 ( .A(n71), .B(n72), .Y(n74) );
  CLKINVX1 U15 ( .A(n118), .Y(n10) );
  CLKINVX1 U16 ( .A(n115), .Y(n4) );
  CLKINVX1 U17 ( .A(n112), .Y(n8) );
  OAI21X1 U18 ( .A0(n11), .A1(n13), .B0(n9), .Y(n112) );
  AOI22X1 U19 ( .A0(n14), .A1(n111), .B0(n13), .B1(n113), .Y(n93) );
  OAI211X1 U21 ( .A0(n15), .A1(n115), .B0(n93), .C0(n3), .Y(n94) );
  CLKINVX1 U22 ( .A(n85), .Y(n14) );
  NAND2X1 U23 ( .A(n97), .B(n6), .Y(n105) );
  NAND2X1 U24 ( .A(n113), .B(n10), .Y(n98) );
  NAND2X1 U25 ( .A(n11), .B(n97), .Y(n107) );
  NAND2X1 U26 ( .A(n118), .B(n85), .Y(n110) );
  OAI21XL U27 ( .A0(n4), .A1(n72), .B0(n108), .Y(n95) );
  CLKINVX1 U28 ( .A(n84), .Y(n7) );
  CLKINVX1 U29 ( .A(addr[2]), .Y(n9) );
  OAI31X1 U30 ( .A0(n71), .A1(addr[6]), .A2(n72), .B0(n87), .Y(n88) );
  OAI21XL U31 ( .A0(n113), .A1(n16), .B0(n14), .Y(n87) );
  OAI211X1 U32 ( .A0(n76), .A1(n71), .B0(n98), .C0(n3), .Y(n77) );
  AOI222XL U35 ( .A0(addr[5]), .A1(addr[6]), .B0(n111), .B1(addr[1]), .C0(n13), 
        .C1(n2), .Y(n76) );
  NAND3XL U36 ( .A(n14), .B(n6), .C(addr[4]), .Y(n117) );
  OAI22XL U37 ( .A0(n116), .A1(n115), .B0(n1), .B1(n112), .Y(n78) );
  CLKINVX3 U38 ( .A(addr[4]), .Y(n71) );
  OAI2BB2XL U39 ( .B0(n115), .B1(n106), .A0N(n72), .A1N(n86), .Y(n89) );
  OAI221XL U40 ( .A0(n116), .A1(addr[4]), .B0(n108), .B1(addr[1]), .C0(n117), 
        .Y(n86) );
  CLKINVX1 U41 ( .A(addr[6]), .Y(n12) );
  CLKINVX1 U42 ( .A(n81), .Y(n5) );
  OAI21XL U44 ( .A0(n96), .A1(n118), .B0(n93), .Y(n82) );
  NAND3X1 U46 ( .A(n101), .B(n100), .C(n99), .Y(n102) );
  AOI32X1 U47 ( .A0(n96), .A1(n6), .A2(n11), .B0(n14), .B1(n95), .Y(n101) );
  AOI2BB2XL U48 ( .B0(n15), .B1(n121), .A0N(n98), .A1N(addr[5]), .Y(n99) );
  OAI21XL U49 ( .A0(n97), .A1(n16), .B0(n13), .Y(n100) );
  AOI2BB2XL U50 ( .B0(n13), .B1(n123), .A0N(n122), .A1N(n9), .Y(n124) );
  AOI211XL U59 ( .A0(n13), .A1(n121), .B0(n120), .C0(n119), .Y(n122) );
  OAI22XL U60 ( .A0(n116), .A1(n115), .B0(addr[5]), .B1(n114), .Y(n120) );
  CLKINVX1 U61 ( .A(n75), .Y(n3) );
  AOI32XL U62 ( .A0(n11), .A1(n96), .A2(n1), .B0(addr[1]), .B1(n121), .Y(n81)
         );
  AOI222XL U63 ( .A0(n13), .A1(n16), .B0(n121), .B1(n116), .C0(n2), .C1(n73), 
        .Y(n80) );
  AOI22XL U64 ( .A0(n78), .A1(n72), .B0(addr[2]), .B1(n77), .Y(n79) );
  NAND2XL U65 ( .A(n111), .B(addr[4]), .Y(n91) );
  AOI211X1 U66 ( .A0(n7), .A1(n110), .B0(n89), .C0(n88), .Y(n90) );
  OAI211X1 U67 ( .A0(n106), .A1(n105), .B0(n104), .C0(n103), .Y(dout[3]) );
  AOI32X1 U68 ( .A0(n2), .A1(n16), .A2(n11), .B0(n94), .B1(n9), .Y(n104) );
  AOI22XL U69 ( .A0(addr[2]), .A1(n102), .B0(n10), .B1(n123), .Y(n103) );
  OAI211X1 U70 ( .A0(addr[2]), .A1(n126), .B0(n125), .C0(n124), .Y(dout[4]) );
  AOI32X1 U71 ( .A0(n14), .A1(n16), .A2(n2), .B0(n8), .B1(n7), .Y(n125) );
  AOI221XL U72 ( .A0(n10), .A1(n111), .B0(n4), .B1(n110), .C0(n109), .Y(n126)
         );
  CLKINVX3 U73 ( .A(n2), .Y(n6) );
  CLKINVX3 U74 ( .A(n106), .Y(n13) );
  CLKINVX3 U75 ( .A(addr[1]), .Y(n15) );
  CLKINVX3 U76 ( .A(n96), .Y(n16) );
endmodule


module sbox5_10 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121;

  OAI222X4 U18 ( .A0(addr[3]), .A1(n106), .B0(n8), .B1(n90), .C0(n13), .C1(n70), .Y(n93) );
  OAI22X2 U40 ( .A0(addr[5]), .A1(n106), .B0(n16), .B1(n114), .Y(n116) );
  NOR2X2 U41 ( .A(n3), .B(addr[3]), .Y(n102) );
  NAND2X2 U45 ( .A(addr[6]), .B(n70), .Y(n114) );
  NAND2X2 U50 ( .A(n70), .B(n8), .Y(n110) );
  NAND2X2 U52 ( .A(addr[1]), .B(n8), .Y(n113) );
  NAND2X2 U54 ( .A(addr[1]), .B(addr[6]), .Y(n106) );
  NAND2X2 U55 ( .A(addr[3]), .B(n13), .Y(n121) );
  CLKINVX1 U1 ( .A(addr[5]), .Y(n1) );
  AOI221XL U2 ( .A0(n93), .A1(n1), .B0(n9), .B1(n14), .C0(n92), .Y(n105) );
  INVX3 U3 ( .A(addr[5]), .Y(n16) );
  OAI221X4 U4 ( .A0(n111), .A1(n110), .B0(n121), .B1(n114), .C0(n109), .Y(n112) );
  OAI221X4 U5 ( .A0(n13), .A1(n114), .B0(n16), .B1(n113), .C0(n120), .Y(n115)
         );
  OAI221X4 U6 ( .A0(n107), .A1(n121), .B0(n111), .B1(n113), .C0(n85), .Y(n86)
         );
  OAI31X1 U7 ( .A0(n68), .A1(addr[5]), .A2(addr[1]), .B0(n81), .Y(n73) );
  OAI32X1 U8 ( .A0(n114), .A1(addr[5]), .A2(n3), .B0(n12), .B1(n107), .Y(n79)
         );
  AOI32XL U9 ( .A0(n14), .A1(n98), .A2(n7), .B0(n2), .B1(n73), .Y(n77) );
  CLKBUFX3 U10 ( .A(addr[4]), .Y(n2) );
  CLKINVX1 U11 ( .A(n81), .Y(n10) );
  NAND2X1 U12 ( .A(n11), .B(n14), .Y(n81) );
  CLKINVX1 U13 ( .A(n110), .Y(n5) );
  CLKXOR2X2 U14 ( .A(n68), .B(n16), .Y(n94) );
  AOI2BB1X1 U15 ( .A0N(n13), .A1N(n1), .B0(n14), .Y(n111) );
  NOR2X1 U16 ( .A(n121), .B(n16), .Y(n91) );
  NOR2BX1 U17 ( .AN(n116), .B(n90), .Y(n83) );
  NAND2X1 U19 ( .A(n5), .B(n16), .Y(n120) );
  CLKINVX1 U20 ( .A(n113), .Y(n7) );
  NAND2X1 U21 ( .A(n7), .B(n16), .Y(n107) );
  CLKINVX1 U22 ( .A(n121), .Y(n12) );
  OAI31X1 U23 ( .A0(n69), .A1(n14), .A2(n113), .B0(n99), .Y(n72) );
  CLKINVX1 U24 ( .A(n106), .Y(n9) );
  OAI2BB2XL U25 ( .B0(n1), .B1(n113), .A0N(n98), .A1N(n11), .Y(n101) );
  CLKINVX1 U26 ( .A(n114), .Y(n11) );
  CLKINVX1 U27 ( .A(n90), .Y(n15) );
  CLKINVX1 U28 ( .A(addr[1]), .Y(n70) );
  CLKINVX1 U29 ( .A(addr[3]), .Y(n68) );
  CLKINVX1 U30 ( .A(addr[6]), .Y(n8) );
  AOI211X1 U31 ( .A0(n91), .A1(addr[1]), .B0(n80), .C0(n79), .Y(n89) );
  OAI2BB2XL U32 ( .B0(n111), .B1(n106), .A0N(n94), .A1N(n5), .Y(n80) );
  AOI211X1 U33 ( .A0(n102), .A1(n84), .B0(n83), .C0(n82), .Y(n85) );
  OAI21XL U34 ( .A0(n8), .A1(n1), .B0(n106), .Y(n84) );
  NOR3XL U35 ( .A(n94), .B(n3), .C(n110), .Y(n82) );
  AOI222XL U36 ( .A0(n9), .A1(n15), .B0(addr[5]), .B1(n108), .C0(n6), .C1(n13), 
        .Y(n109) );
  CLKINVX1 U37 ( .A(n107), .Y(n6) );
  OAI21XL U38 ( .A0(addr[6]), .A1(addr[3]), .B0(n106), .Y(n108) );
  NAND2X1 U39 ( .A(addr[3]), .B(n3), .Y(n90) );
  NAND2X1 U42 ( .A(n2), .B(addr[5]), .Y(n98) );
  NAND2X1 U43 ( .A(n3), .B(n68), .Y(n97) );
  OAI21XL U44 ( .A0(addr[1]), .A1(n97), .B0(n96), .Y(n103) );
  AOI33XL U46 ( .A0(n3), .A1(n95), .A2(addr[5]), .B0(n94), .B1(n13), .B2(
        addr[1]), .Y(n96) );
  OAI21XL U47 ( .A0(n70), .A1(n68), .B0(n114), .Y(n95) );
  OAI21XL U48 ( .A0(addr[6]), .A1(n121), .B0(n99), .Y(n100) );
  NAND2X1 U49 ( .A(n71), .B(n5), .Y(n99) );
  XOR2X1 U51 ( .A(n69), .B(n3), .Y(n71) );
  AOI2BB2XL U53 ( .B0(n102), .B1(n116), .A0N(n2), .A1N(n75), .Y(n76) );
  AOI211X1 U56 ( .A0(n4), .A1(n3), .B0(n74), .C0(n83), .Y(n75) );
  AO22XL U57 ( .A0(n7), .A1(n12), .B0(addr[6]), .B1(n102), .Y(n74) );
  CLKINVX1 U58 ( .A(n120), .Y(n4) );
  CLKINVX1 U59 ( .A(n2), .Y(n69) );
  AO22XL U60 ( .A0(n7), .A1(n15), .B0(addr[6]), .B1(n91), .Y(n92) );
  AOI222XL U61 ( .A0(n116), .A1(n13), .B0(addr[3]), .B1(n115), .C0(n7), .C1(
        n14), .Y(n117) );
  OAI221X1 U62 ( .A0(n2), .A1(n105), .B0(n110), .B1(n121), .C0(n104), .Y(
        dout[3]) );
  AOI222XL U63 ( .A0(n2), .A1(n103), .B0(n102), .B1(n101), .C0(n100), .C1(n1), 
        .Y(n104) );
  OAI211X1 U64 ( .A0(n2), .A1(n89), .B0(n88), .C0(n87), .Y(dout[2]) );
  AOI33XL U65 ( .A0(n12), .A1(n98), .A2(n11), .B0(n3), .B1(n94), .B2(n5), .Y(
        n88) );
  AOI222XL U66 ( .A0(n10), .A1(n16), .B0(n2), .B1(n86), .C0(n91), .C1(n9), .Y(
        n87) );
  OAI211X1 U67 ( .A0(n78), .A1(n16), .B0(n77), .C0(n76), .Y(dout[1]) );
  AOI221XL U68 ( .A0(n12), .A1(addr[1]), .B0(n9), .B1(n14), .C0(n72), .Y(n78)
         );
  OAI211X1 U69 ( .A0(n121), .A1(n120), .B0(n119), .C0(n118), .Y(dout[4]) );
  AOI32XL U70 ( .A0(n14), .A1(n114), .A2(addr[5]), .B0(n2), .B1(n112), .Y(n119) );
  AOI2BB2X1 U71 ( .B0(n10), .B1(n16), .A0N(n2), .A1N(n117), .Y(n118) );
  BUFX4 U72 ( .A(addr[2]), .Y(n3) );
  CLKINVX3 U73 ( .A(n3), .Y(n13) );
  CLKINVX3 U74 ( .A(n97), .Y(n14) );
endmodule


module sbox6_10 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147;

  NAND2X2 U39 ( .A(n138), .B(addr[3]), .Y(n147) );
  NOR2X2 U47 ( .A(n7), .B(n17), .Y(n138) );
  NOR2X2 U50 ( .A(n13), .B(n4), .Y(n119) );
  NOR2X2 U58 ( .A(n84), .B(n13), .Y(n125) );
  NAND2X2 U61 ( .A(n97), .B(n103), .Y(n112) );
  NOR2X2 U62 ( .A(n85), .B(addr[1]), .Y(n103) );
  NOR2X2 U63 ( .A(n84), .B(addr[3]), .Y(n97) );
  NAND2X2 U64 ( .A(n117), .B(n131), .Y(n140) );
  NOR2X2 U65 ( .A(n5), .B(addr[3]), .Y(n131) );
  NOR2X2 U66 ( .A(n18), .B(addr[6]), .Y(n117) );
  NOR2X1 U1 ( .A(n7), .B(addr[3]), .Y(n102) );
  AOI211X1 U2 ( .A0(n15), .A1(n13), .B0(n131), .C0(n143), .Y(n121) );
  CLKINVX1 U3 ( .A(addr[3]), .Y(n1) );
  INVX3 U4 ( .A(addr[3]), .Y(n13) );
  CLKINVX1 U5 ( .A(n84), .Y(n2) );
  INVX4 U6 ( .A(n4), .Y(n84) );
  CLKBUFX3 U7 ( .A(addr[4]), .Y(n4) );
  CLKINVX1 U8 ( .A(n7), .Y(n3) );
  OAI222X1 U9 ( .A0(n91), .A1(n15), .B0(n5), .B1(n14), .C0(addr[5]), .C1(n11), 
        .Y(n92) );
  BUFX4 U10 ( .A(addr[2]), .Y(n5) );
  OAI221X1 U11 ( .A0(n85), .A1(n12), .B0(n13), .B1(n16), .C0(n86), .Y(n90) );
  INVX3 U12 ( .A(n96), .Y(n16) );
  OAI221X4 U13 ( .A0(n123), .A1(n82), .B0(n17), .B1(n15), .C0(n9), .Y(n124) );
  NOR2X4 U14 ( .A(addr[1]), .B(addr[6]), .Y(n130) );
  NOR2X4 U15 ( .A(n5), .B(addr[5]), .Y(n143) );
  INVX1 U16 ( .A(n130), .Y(n83) );
  CLKINVX1 U17 ( .A(n125), .Y(n12) );
  NAND2X1 U18 ( .A(n83), .B(n16), .Y(n105) );
  INVXL U19 ( .A(n121), .Y(n8) );
  CLKINVX1 U20 ( .A(n138), .Y(n6) );
  CLKINVX1 U21 ( .A(n117), .Y(n17) );
  CLKINVX1 U22 ( .A(n119), .Y(n11) );
  NOR2X1 U23 ( .A(n16), .B(n123), .Y(n144) );
  NOR2X1 U24 ( .A(n18), .B(n85), .Y(n96) );
  CLKINVX1 U25 ( .A(n103), .Y(n82) );
  OAI211X1 U26 ( .A0(n83), .A1(n12), .B0(n104), .C0(n112), .Y(n108) );
  OAI21XL U27 ( .A0(n103), .A1(n117), .B0(n102), .Y(n104) );
  OAI21XL U28 ( .A0(n132), .A1(n85), .B0(n1), .Y(n86) );
  AOI21X1 U29 ( .A0(n84), .A1(n102), .B0(n125), .Y(n91) );
  OAI2BB2XL U30 ( .B0(n143), .B1(n83), .A0N(n143), .A1N(n117), .Y(n118) );
  CLKINVX1 U31 ( .A(n122), .Y(n9) );
  CLKINVX1 U32 ( .A(n126), .Y(n81) );
  CLKINVX1 U33 ( .A(n97), .Y(n14) );
  NAND2BX1 U34 ( .AN(n144), .B(n137), .Y(n107) );
  CLKINVX1 U35 ( .A(addr[1]), .Y(n18) );
  NOR2X1 U36 ( .A(n16), .B(n3), .Y(n122) );
  NOR2X1 U37 ( .A(addr[1]), .B(n2), .Y(n132) );
  OAI22X1 U38 ( .A0(n11), .A1(n17), .B0(n5), .B1(n81), .Y(n88) );
  NAND2X1 U40 ( .A(n3), .B(n15), .Y(n123) );
  NAND4X1 U41 ( .A(n147), .B(n140), .C(n100), .D(n99), .Y(n101) );
  AOI222XL U42 ( .A0(n98), .A1(n7), .B0(n102), .B1(n130), .C0(n97), .C1(n105), 
        .Y(n99) );
  NAND3X1 U43 ( .A(n5), .B(n11), .C(n96), .Y(n100) );
  OAI221X1 U44 ( .A0(n13), .A1(n82), .B0(n11), .B1(n85), .C0(n81), .Y(n98) );
  AOI22X1 U45 ( .A0(n4), .A1(n115), .B0(addr[5]), .B1(n114), .Y(n129) );
  OAI21XL U46 ( .A0(n121), .A1(n83), .B0(n147), .Y(n115) );
  OAI21XL U48 ( .A0(n113), .A1(n7), .B0(n112), .Y(n114) );
  AOI221XL U49 ( .A0(n119), .A1(n18), .B0(n130), .B1(addr[3]), .C0(n111), .Y(
        n113) );
  OAI22XL U51 ( .A0(n17), .A1(n84), .B0(addr[3]), .B1(n16), .Y(n111) );
  OAI22XL U52 ( .A0(n13), .A1(n85), .B0(addr[1]), .B1(n11), .Y(n142) );
  AOI211X1 U53 ( .A0(n4), .A1(n135), .B0(n134), .C0(n133), .Y(n136) );
  OA21XL U54 ( .A0(n1), .A1(n3), .B0(n132), .Y(n133) );
  OAI2BB2XL U55 ( .B0(n2), .B1(n9), .A0N(n131), .A1N(n130), .Y(n134) );
  OAI22X1 U56 ( .A0(n5), .A1(n17), .B0(n7), .B1(n16), .Y(n135) );
  CLKINVX3 U57 ( .A(addr[5]), .Y(n15) );
  AOI2BB2X1 U59 ( .B0(n5), .B1(n130), .A0N(n3), .A1N(n82), .Y(n137) );
  NOR2X1 U60 ( .A(n82), .B(n2), .Y(n126) );
  AOI2BB2XL U67 ( .B0(n143), .B1(n90), .A0N(n89), .A1N(n15), .Y(n94) );
  AOI211X1 U68 ( .A0(n122), .A1(n4), .B0(n88), .C0(n87), .Y(n89) );
  OAI32X1 U69 ( .A0(n82), .A1(n13), .A2(n7), .B0(n6), .B1(n14), .Y(n87) );
  NAND3X1 U70 ( .A(n147), .B(n140), .C(n139), .Y(n141) );
  AOI32X1 U71 ( .A0(n5), .A1(n18), .A2(n4), .B0(n138), .B1(n84), .Y(n139) );
  AO22XL U72 ( .A0(n143), .A1(n2), .B0(n116), .B1(n84), .Y(n120) );
  OAI21XL U73 ( .A0(n3), .A1(n15), .B0(n123), .Y(n116) );
  CLKINVX1 U74 ( .A(n106), .Y(n10) );
  AOI32XL U75 ( .A0(n105), .A1(n84), .A2(n1), .B0(addr[1]), .B1(n125), .Y(n106) );
  OAI211X1 U76 ( .A0(n84), .A1(n140), .B0(n110), .C0(n109), .Y(dout[2]) );
  AOI222XL U77 ( .A0(n108), .A1(n15), .B0(n143), .B1(n10), .C0(n119), .C1(n107), .Y(n109) );
  AOI2BB2XL U78 ( .B0(addr[5]), .B1(n101), .A0N(n7), .A1N(n112), .Y(n110) );
  OAI211X1 U79 ( .A0(n2), .A1(n147), .B0(n146), .C0(n145), .Y(dout[4]) );
  AOI222XL U80 ( .A0(n144), .A1(n13), .B0(n143), .B1(n142), .C0(n141), .C1(n15), .Y(n145) );
  OA22X1 U81 ( .A0(n12), .A1(n137), .B0(n136), .B1(n15), .Y(n146) );
  NAND3X1 U82 ( .A(n129), .B(n128), .C(n127), .Y(dout[3]) );
  AOI32XL U83 ( .A0(n120), .A1(n13), .A2(addr[1]), .B0(n119), .B1(n118), .Y(
        n128) );
  AOI222XL U84 ( .A0(n144), .A1(n84), .B0(n126), .B1(n8), .C0(n125), .C1(n124), 
        .Y(n127) );
  NAND3BX1 U85 ( .AN(n95), .B(n94), .C(n93), .Y(dout[1]) );
  OAI222X1 U86 ( .A0(n140), .A1(n4), .B0(n112), .B1(n7), .C0(n16), .C1(n91), 
        .Y(n95) );
  AOI32XL U87 ( .A0(addr[1]), .A1(n15), .A2(n125), .B0(n130), .B1(n92), .Y(n93) );
  CLKINVX3 U88 ( .A(n5), .Y(n7) );
  CLKINVX3 U89 ( .A(addr[6]), .Y(n85) );
endmodule


module sbox7_10 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148;

  OAI222X4 U19 ( .A0(n11), .A1(n129), .B0(n4), .B1(n7), .C0(addr[1]), .C1(n18), 
        .Y(n122) );
  OAI33X4 U33 ( .A0(addr[1]), .A1(n4), .A2(n5), .B0(n8), .B1(n86), .B2(n12), 
        .Y(n97) );
  NOR2X2 U44 ( .A(n16), .B(n4), .Y(n116) );
  NOR2X2 U48 ( .A(addr[1]), .B(addr[6]), .Y(n136) );
  NOR2X2 U51 ( .A(n21), .B(n16), .Y(n125) );
  NOR2X2 U52 ( .A(n8), .B(addr[3]), .Y(n131) );
  NOR2X2 U58 ( .A(n93), .B(n124), .Y(n142) );
  NOR2X2 U60 ( .A(n85), .B(addr[1]), .Y(n93) );
  NOR2X2 U62 ( .A(n87), .B(n3), .Y(n137) );
  NOR2X2 U65 ( .A(n85), .B(n9), .Y(n140) );
  NAND2X1 U1 ( .A(n3), .B(n4), .Y(n119) );
  CLKBUFX3 U2 ( .A(addr[4]), .Y(n4) );
  CLKINVX1 U3 ( .A(n87), .Y(n1) );
  CLKINVX1 U4 ( .A(n86), .Y(n2) );
  CLKBUFX3 U5 ( .A(addr[2]), .Y(n5) );
  OAI31X1 U6 ( .A0(n16), .A1(n87), .A2(n9), .B0(n117), .Y(n121) );
  OAI22X1 U7 ( .A0(addr[1]), .A1(n18), .B0(n5), .B1(n113), .Y(n100) );
  OAI22X1 U8 ( .A0(n4), .A1(n21), .B0(addr[3]), .B1(n84), .Y(n103) );
  NOR2X4 U9 ( .A(n9), .B(addr[6]), .Y(n124) );
  AOI211XL U10 ( .A0(n5), .A1(n6), .B0(n131), .C0(n130), .Y(n132) );
  NOR3XL U11 ( .A(n11), .B(addr[3]), .C(n2), .Y(n130) );
  OAI21XL U12 ( .A0(n3), .A1(n1), .B0(n119), .Y(n89) );
  BUFX4 U13 ( .A(addr[5]), .Y(n3) );
  AOI221XL U14 ( .A0(n140), .A1(n89), .B0(n109), .B1(n6), .C0(n88), .Y(n96) );
  CLKINVX1 U15 ( .A(n140), .Y(n8) );
  OAI2BB2XL U16 ( .B0(n142), .B1(n84), .A0N(n141), .A1N(n140), .Y(n143) );
  CLKINVX1 U17 ( .A(n125), .Y(n14) );
  CLKINVX1 U18 ( .A(n142), .Y(n6) );
  NAND2X1 U20 ( .A(n14), .B(n19), .Y(n105) );
  CLKINVX1 U21 ( .A(n123), .Y(n17) );
  CLKINVX1 U22 ( .A(n109), .Y(n15) );
  NAND2X1 U23 ( .A(n124), .B(n16), .Y(n113) );
  CLKINVX1 U24 ( .A(n137), .Y(n84) );
  NOR2X1 U25 ( .A(n84), .B(n16), .Y(n109) );
  CLKINVX1 U26 ( .A(n136), .Y(n11) );
  OAI22XL U27 ( .A0(n137), .A1(n7), .B0(n9), .B1(n15), .Y(n146) );
  OAI21X1 U28 ( .A0(n87), .A1(n14), .B0(n129), .Y(n141) );
  NAND2X1 U29 ( .A(n116), .B(n21), .Y(n129) );
  CLKINVX1 U30 ( .A(n93), .Y(n10) );
  OAI21XL U31 ( .A0(n119), .A1(n10), .B0(n118), .Y(n120) );
  OAI21XL U32 ( .A0(n125), .A1(n137), .B0(n124), .Y(n118) );
  NOR2X1 U34 ( .A(n21), .B(n18), .Y(n123) );
  CLKINVX1 U35 ( .A(n145), .Y(n18) );
  OAI22XL U36 ( .A0(n137), .A1(n113), .B0(n85), .B1(n17), .Y(n88) );
  CLKINVX1 U37 ( .A(n116), .Y(n12) );
  CLKINVX1 U38 ( .A(n131), .Y(n7) );
  CLKINVX1 U39 ( .A(n134), .Y(n19) );
  NOR2XL U40 ( .A(n125), .B(n87), .Y(n110) );
  CLKINVX1 U41 ( .A(n119), .Y(n83) );
  CLKINVX1 U42 ( .A(n103), .Y(n20) );
  OA21XL U43 ( .A0(n13), .A1(n10), .B0(n117), .Y(n102) );
  CLKINVX1 U45 ( .A(n105), .Y(n13) );
  OAI2BB1XL U46 ( .A0N(n103), .A1N(n124), .B0(n102), .Y(n104) );
  OAI22X1 U47 ( .A0(n21), .A1(n12), .B0(n4), .B1(n19), .Y(n112) );
  NOR4X1 U49 ( .A(n4), .B(addr[3]), .C(n9), .D(n86), .Y(n99) );
  XNOR2X1 U50 ( .A(addr[6]), .B(n5), .Y(n101) );
  AOI211X1 U53 ( .A0(n116), .A1(addr[6]), .B0(n115), .C0(n114), .Y(n128) );
  OAI222X1 U54 ( .A0(n111), .A1(n8), .B0(n110), .B1(n10), .C0(n11), .C1(n15), 
        .Y(n115) );
  OAI2BB2XL U55 ( .B0(n83), .B1(n113), .A0N(n9), .A1N(n112), .Y(n114) );
  OA21XL U56 ( .A0(n16), .A1(n3), .B0(n17), .Y(n111) );
  NAND2X1 U57 ( .A(n5), .B(n136), .Y(n133) );
  CLKINVX1 U59 ( .A(addr[6]), .Y(n85) );
  AOI211X1 U61 ( .A0(n131), .A1(n3), .B0(n92), .C0(n91), .Y(n95) );
  OAI221X1 U63 ( .A0(n9), .A1(n18), .B0(n8), .B1(n84), .C0(n102), .Y(n92) );
  OAI31X1 U64 ( .A0(n16), .A1(n87), .A2(n11), .B0(n90), .Y(n91) );
  AO21XL U66 ( .A0(n119), .A1(n129), .B0(addr[6]), .Y(n90) );
  NOR2X1 U67 ( .A(n87), .B(addr[3]), .Y(n145) );
  AOI21XL U68 ( .A0(addr[3]), .A1(n98), .B0(n97), .Y(n108) );
  OAI2BB1XL U69 ( .A0N(n86), .A1N(n124), .B0(n133), .Y(n98) );
  NAND3X1 U70 ( .A(n136), .B(n16), .C(n3), .Y(n117) );
  NOR2X1 U71 ( .A(addr[3]), .B(n3), .Y(n134) );
  OAI21X1 U72 ( .A0(n5), .A1(n142), .B0(n133), .Y(n138) );
  OAI22XL U73 ( .A0(n142), .A1(n12), .B0(n1), .B1(n132), .Y(n135) );
  AO21X1 U74 ( .A0(n139), .A1(n21), .B0(n138), .Y(n144) );
  OAI21XL U75 ( .A0(n2), .A1(n9), .B0(n10), .Y(n139) );
  OAI221X1 U76 ( .A0(n96), .A1(n86), .B0(n5), .B1(n95), .C0(n94), .Y(dout[1])
         );
  AOI2BB2X1 U77 ( .B0(n93), .B1(n112), .A0N(n133), .A1N(n20), .Y(n94) );
  OAI211X1 U78 ( .A0(n128), .A1(n86), .B0(n127), .C0(n126), .Y(dout[3]) );
  AOI32XL U79 ( .A0(n125), .A1(n1), .A2(n124), .B0(n123), .B1(n136), .Y(n126)
         );
  OAI31X1 U80 ( .A0(n122), .A1(n121), .A2(n120), .B0(n86), .Y(n127) );
  OAI221X1 U81 ( .A0(n3), .A1(n108), .B0(n107), .B1(n21), .C0(n106), .Y(
        dout[2]) );
  AOI32XL U82 ( .A0(n105), .A1(n86), .A2(n140), .B0(n2), .B1(n104), .Y(n106)
         );
  AOI211X1 U83 ( .A0(n101), .A1(n4), .B0(n100), .C0(n99), .Y(n107) );
  NAND2X1 U84 ( .A(n148), .B(n147), .Y(dout[4]) );
  AOI222XL U85 ( .A0(n136), .A1(n141), .B0(n3), .B1(n135), .C0(n134), .C1(n138), .Y(n148) );
  AOI222XL U86 ( .A0(n5), .A1(n146), .B0(n145), .B1(n144), .C0(n143), .C1(n86), 
        .Y(n147) );
  CLKINVX3 U87 ( .A(addr[1]), .Y(n9) );
  CLKINVX3 U88 ( .A(addr[3]), .Y(n16) );
  CLKINVX3 U89 ( .A(n3), .Y(n21) );
  CLKINVX3 U90 ( .A(n5), .Y(n86) );
  CLKINVX3 U91 ( .A(n4), .Y(n87) );
endmodule


module sbox8_10 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132;

  NAND2X2 U41 ( .A(addr[6]), .B(n10), .Y(n131) );
  NAND2X2 U48 ( .A(addr[4]), .B(n16), .Y(n123) );
  NAND2X2 U49 ( .A(n2), .B(n74), .Y(n87) );
  NAND2X2 U50 ( .A(addr[1]), .B(n6), .Y(n124) );
  NAND2X2 U54 ( .A(addr[2]), .B(n75), .Y(n116) );
  NAND2X2 U60 ( .A(addr[6]), .B(addr[1]), .Y(n105) );
  NAND2X2 U61 ( .A(n10), .B(n6), .Y(n108) );
  OAI31X1 U1 ( .A0(n123), .A1(addr[6]), .A2(n116), .B0(n109), .Y(n110) );
  AOI222X1 U2 ( .A0(n88), .A1(addr[2]), .B0(n74), .B1(n11), .C0(n12), .C1(n92), 
        .Y(n114) );
  OAI222X1 U3 ( .A0(addr[2]), .A1(n126), .B0(n16), .B1(n125), .C0(n124), .C1(
        n123), .Y(n127) );
  NAND2X4 U4 ( .A(addr[4]), .B(n2), .Y(n115) );
  OAI32X1 U5 ( .A0(n6), .A1(addr[4]), .A2(n92), .B0(n115), .B1(n108), .Y(n96)
         );
  OAI221X1 U6 ( .A0(n105), .A1(n87), .B0(addr[4]), .B1(n108), .C0(n86), .Y(n90) );
  AOI32XL U7 ( .A0(n4), .A1(n14), .A2(n2), .B0(n5), .B1(n117), .Y(n130) );
  OA21XL U8 ( .A0(n12), .A1(n75), .B0(n121), .Y(n78) );
  INVXL U9 ( .A(n119), .Y(n3) );
  INVX3 U10 ( .A(n2), .Y(n16) );
  BUFX4 U11 ( .A(addr[3]), .Y(n2) );
  CLKBUFX3 U12 ( .A(addr[5]), .Y(n1) );
  CLKINVX1 U13 ( .A(n108), .Y(n5) );
  CLKINVX1 U14 ( .A(n107), .Y(n13) );
  CLKINVX1 U15 ( .A(n93), .Y(n15) );
  NAND2X1 U16 ( .A(n16), .B(n74), .Y(n93) );
  NAND2X1 U17 ( .A(n12), .B(n75), .Y(n121) );
  OAI21XL U18 ( .A0(n115), .A1(n75), .B0(n107), .Y(n77) );
  OAI21X1 U19 ( .A0(n74), .A1(n75), .B0(n123), .Y(n88) );
  OAI31XL U20 ( .A0(n115), .A1(n10), .A2(n116), .B0(n118), .Y(n94) );
  CLKINVX1 U21 ( .A(n131), .Y(n9) );
  NAND2X1 U22 ( .A(n14), .B(n16), .Y(n107) );
  OAI22XL U23 ( .A0(n116), .A1(n123), .B0(n14), .B1(n115), .Y(n117) );
  OAI22XL U24 ( .A0(n123), .A1(n108), .B0(n131), .B1(n93), .Y(n95) );
  OAI2BB2XL U25 ( .B0(n115), .B1(n131), .A0N(n88), .A1N(n8), .Y(n89) );
  AOI211XL U26 ( .A0(n108), .A1(n105), .B0(n74), .C0(n121), .Y(n85) );
  CLKINVX1 U27 ( .A(n124), .Y(n4) );
  OAI22XL U28 ( .A0(n14), .A1(n123), .B0(n78), .B1(n87), .Y(n81) );
  NAND2BX2 U29 ( .AN(n78), .B(n16), .Y(n120) );
  NAND2XL U30 ( .A(n115), .B(n93), .Y(n104) );
  OAI2BB2XL U31 ( .B0(n106), .B1(n105), .A0N(n104), .A1N(n4), .Y(n111) );
  NOR2BXL U32 ( .AN(n123), .B(n103), .Y(n106) );
  NAND3X1 U33 ( .A(n104), .B(n10), .C(n14), .Y(n84) );
  AO21X1 U34 ( .A0(n14), .A1(n8), .B0(n101), .Y(n102) );
  OAI33X1 U35 ( .A0(n6), .A1(n16), .A2(n100), .B0(n12), .B1(n103), .B2(n124), 
        .Y(n101) );
  OA22XL U36 ( .A0(n107), .A1(n131), .B0(n120), .B1(n124), .Y(n98) );
  CLKINVX1 U37 ( .A(n125), .Y(n7) );
  OAI21XL U38 ( .A0(n4), .A1(n9), .B0(addr[4]), .Y(n86) );
  NAND2X1 U39 ( .A(n1), .B(n12), .Y(n100) );
  OAI221X1 U40 ( .A0(n124), .A1(n121), .B0(addr[1]), .B1(n120), .C0(n3), .Y(
        n128) );
  OAI31XL U42 ( .A0(n12), .A1(n10), .A2(n16), .B0(n118), .Y(n119) );
  NAND2X1 U43 ( .A(n8), .B(addr[2]), .Y(n125) );
  NAND4XL U44 ( .A(n9), .B(n1), .C(n2), .D(addr[2]), .Y(n109) );
  NAND3X1 U45 ( .A(n14), .B(n6), .C(n2), .Y(n118) );
  OAI21XL U46 ( .A0(n1), .A1(n87), .B0(n114), .Y(n76) );
  OAI22XL U47 ( .A0(n108), .A1(n120), .B0(n79), .B1(n100), .Y(n80) );
  AOI221XL U51 ( .A0(n9), .A1(n16), .B0(n8), .B1(n2), .C0(n91), .Y(n79) );
  NOR2X1 U52 ( .A(n1), .B(n2), .Y(n103) );
  NOR2X1 U53 ( .A(n87), .B(addr[6]), .Y(n91) );
  NOR2X1 U55 ( .A(n16), .B(n1), .Y(n92) );
  CLKINVX1 U56 ( .A(n100), .Y(n11) );
  OA21XL U57 ( .A0(n1), .A1(n115), .B0(n120), .Y(n132) );
  AOI221XL U58 ( .A0(n5), .A1(n2), .B0(n8), .B1(addr[4]), .C0(n122), .Y(n126)
         );
  OAI22XL U59 ( .A0(n2), .A1(n10), .B0(addr[4]), .B1(n131), .Y(n122) );
  OAI211X1 U62 ( .A0(addr[2]), .A1(n99), .B0(n98), .C0(n97), .Y(dout[2]) );
  AOI221XL U63 ( .A0(addr[2]), .A1(n96), .B0(n1), .B1(n95), .C0(n94), .Y(n97)
         );
  AOI221XL U64 ( .A0(n91), .A1(n1), .B0(n90), .B1(n75), .C0(n89), .Y(n99) );
  OAI211X1 U65 ( .A0(n132), .A1(n131), .B0(n130), .C0(n129), .Y(dout[4]) );
  AOI222XL U66 ( .A0(n128), .A1(n74), .B0(n1), .B1(n127), .C0(n13), .C1(n8), 
        .Y(n129) );
  OAI211X1 U67 ( .A0(addr[1]), .A1(n114), .B0(n113), .C0(n112), .Y(dout[3]) );
  AOI221XL U68 ( .A0(n111), .A1(n12), .B0(n13), .B1(n5), .C0(n110), .Y(n112)
         );
  AOI2BB2XL U69 ( .B0(n102), .B1(n74), .A0N(n115), .A1N(n125), .Y(n113) );
  NAND4BX1 U70 ( .AN(n85), .B(n84), .C(n83), .D(n82), .Y(dout[1]) );
  AOI221XL U71 ( .A0(n9), .A1(n81), .B0(n15), .B1(n7), .C0(n80), .Y(n82) );
  AOI22X1 U72 ( .A0(n8), .A1(n77), .B0(n4), .B1(n76), .Y(n83) );
  CLKINVX3 U73 ( .A(addr[6]), .Y(n6) );
  CLKINVX3 U74 ( .A(n105), .Y(n8) );
  CLKINVX3 U75 ( .A(addr[1]), .Y(n10) );
  CLKINVX3 U76 ( .A(addr[2]), .Y(n12) );
  CLKINVX3 U77 ( .A(n116), .Y(n14) );
  CLKINVX3 U78 ( .A(addr[4]), .Y(n74) );
  CLKINVX3 U79 ( .A(n1), .Y(n75) );
endmodule


module crp_10 ( P, R, K_sub );
  output [1:32] P;
  input [1:32] R;
  input [1:48] K_sub;
  wire   n1;
  wire   [1:48] X;

  sbox1_10 u0 ( .addr(X[1:6]), .dout({P[9], P[17], P[23], P[31]}) );
  sbox2_10 u1 ( .addr({X[7], n1, X[9:12]}), .dout({P[13], P[28], P[2], P[18]})
         );
  sbox3_10 u2 ( .addr(X[13:18]), .dout({P[24], P[16], P[30], P[6]}) );
  sbox4_10 u3 ( .addr(X[19:24]), .dout({P[26], P[20], P[10], P[1]}) );
  sbox5_10 u4 ( .addr(X[25:30]), .dout({P[8], P[14], P[25], P[3]}) );
  sbox6_10 u5 ( .addr(X[31:36]), .dout({P[4], P[29], P[11], P[19]}) );
  sbox7_10 u6 ( .addr(X[37:42]), .dout({P[32], P[12], P[22], P[7]}) );
  sbox8_10 u7 ( .addr(X[43:48]), .dout({P[5], P[27], P[15], P[21]}) );
  XNOR2X1 U1 ( .A(R[5]), .B(K_sub[8]), .Y(X[8]) );
  INVX3 U2 ( .A(X[8]), .Y(n1) );
  XOR2X1 U3 ( .A(R[1]), .B(K_sub[2]), .Y(X[2]) );
  CLKXOR2X4 U4 ( .A(R[29]), .B(K_sub[42]), .Y(X[42]) );
  CLKXOR2X4 U5 ( .A(R[16]), .B(K_sub[25]), .Y(X[25]) );
  CLKXOR2X4 U6 ( .A(R[8]), .B(K_sub[11]), .Y(X[11]) );
  CLKXOR2X4 U7 ( .A(R[22]), .B(K_sub[33]), .Y(X[33]) );
  CLKXOR2X4 U8 ( .A(R[29]), .B(K_sub[44]), .Y(X[44]) );
  CLKXOR2X4 U9 ( .A(R[16]), .B(K_sub[23]), .Y(X[23]) );
  CLKXOR2X4 U10 ( .A(R[26]), .B(K_sub[39]), .Y(X[39]) );
  CLKXOR2X4 U11 ( .A(R[10]), .B(K_sub[15]), .Y(X[15]) );
  CLKXOR2X4 U12 ( .A(R[20]), .B(K_sub[31]), .Y(X[31]) );
  CLKXOR2X4 U13 ( .A(R[31]), .B(K_sub[46]), .Y(X[46]) );
  CLKXOR2X4 U14 ( .A(R[12]), .B(K_sub[19]), .Y(X[19]) );
  CLKXOR2X4 U15 ( .A(R[20]), .B(K_sub[29]), .Y(X[29]) );
  CLKXOR2X2 U16 ( .A(R[4]), .B(K_sub[5]), .Y(X[5]) );
  CLKXOR2X2 U17 ( .A(R[15]), .B(K_sub[22]), .Y(X[22]) );
  CLKXOR2X2 U18 ( .A(R[24]), .B(K_sub[35]), .Y(X[35]) );
  CLKXOR2X2 U19 ( .A(R[21]), .B(K_sub[30]), .Y(X[30]) );
  CLKXOR2X2 U20 ( .A(R[12]), .B(K_sub[17]), .Y(X[17]) );
  CLKXOR2X2 U21 ( .A(R[32]), .B(K_sub[1]), .Y(X[1]) );
  CLKXOR2X2 U22 ( .A(R[13]), .B(K_sub[20]), .Y(X[20]) );
  CLKXOR2X2 U23 ( .A(R[18]), .B(K_sub[27]), .Y(X[27]) );
  CLKXOR2X2 U24 ( .A(R[8]), .B(K_sub[13]), .Y(X[13]) );
  CLKXOR2X2 U25 ( .A(R[5]), .B(K_sub[6]), .Y(X[6]) );
  CLKXOR2X2 U26 ( .A(R[4]), .B(K_sub[7]), .Y(X[7]) );
  CLKXOR2X2 U27 ( .A(R[24]), .B(K_sub[37]), .Y(X[37]) );
  CLKXOR2X2 U28 ( .A(R[28]), .B(K_sub[43]), .Y(X[43]) );
  CLKXOR2X2 U29 ( .A(R[1]), .B(K_sub[48]), .Y(X[48]) );
  CLKXOR2X2 U30 ( .A(R[17]), .B(K_sub[24]), .Y(X[24]) );
  CLKXOR2X2 U31 ( .A(R[9]), .B(K_sub[12]), .Y(X[12]) );
  CLKXOR2X2 U32 ( .A(R[13]), .B(K_sub[18]), .Y(X[18]) );
  CLKXOR2X2 U33 ( .A(R[25]), .B(K_sub[36]), .Y(X[36]) );
  XOR2X1 U34 ( .A(R[23]), .B(K_sub[34]), .Y(X[34]) );
  XOR2X1 U35 ( .A(R[9]), .B(K_sub[14]), .Y(X[14]) );
  XOR2X1 U36 ( .A(R[30]), .B(K_sub[45]), .Y(X[45]) );
  XOR2X1 U37 ( .A(R[21]), .B(K_sub[32]), .Y(X[32]) );
  XOR2X1 U38 ( .A(R[25]), .B(K_sub[38]), .Y(X[38]) );
  XOR2X1 U39 ( .A(R[27]), .B(K_sub[40]), .Y(X[40]) );
  XOR2X1 U40 ( .A(R[3]), .B(K_sub[4]), .Y(X[4]) );
  XOR2X1 U41 ( .A(R[11]), .B(K_sub[16]), .Y(X[16]) );
  XOR2X1 U42 ( .A(R[7]), .B(K_sub[10]), .Y(X[10]) );
  XOR2X1 U43 ( .A(R[14]), .B(K_sub[21]), .Y(X[21]) );
  XOR2X1 U44 ( .A(R[6]), .B(K_sub[9]), .Y(X[9]) );
  XOR2X1 U45 ( .A(R[2]), .B(K_sub[3]), .Y(X[3]) );
  XOR2X1 U46 ( .A(R[28]), .B(K_sub[41]), .Y(X[41]) );
  XOR2X1 U47 ( .A(R[17]), .B(K_sub[26]), .Y(X[26]) );
  XOR2X1 U48 ( .A(R[32]), .B(K_sub[47]), .Y(X[47]) );
  XOR2X1 U49 ( .A(R[19]), .B(K_sub[28]), .Y(X[28]) );
endmodule


module sbox1_9 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127;

  OAI222X4 U13 ( .A0(addr[5]), .A1(n101), .B0(n1), .B1(n100), .C0(n99), .C1(n8), .Y(dout[3]) );
  OAI21X2 U42 ( .A0(n4), .A1(n112), .B0(n106), .Y(n123) );
  NAND2X2 U44 ( .A(addr[6]), .B(n70), .Y(n115) );
  NAND2X2 U48 ( .A(addr[1]), .B(n11), .Y(n114) );
  OAI22X2 U49 ( .A0(n71), .A1(n6), .B0(addr[5]), .B1(n120), .Y(n85) );
  NAND2X2 U50 ( .A(n3), .B(n71), .Y(n120) );
  NOR2X2 U51 ( .A(n71), .B(n3), .Y(n124) );
  NOR3X2 U55 ( .A(n2), .B(addr[6]), .C(n8), .Y(n102) );
  NOR2X2 U56 ( .A(n109), .B(n3), .Y(n93) );
  NAND2X2 U57 ( .A(addr[1]), .B(addr[6]), .Y(n109) );
  NAND2X2 U59 ( .A(n70), .B(n11), .Y(n112) );
  NOR2X1 U1 ( .A(n114), .B(n120), .Y(n104) );
  BUFX4 U2 ( .A(addr[4]), .Y(n2) );
  CLKBUFX3 U3 ( .A(addr[2]), .Y(n1) );
  OAI32X1 U4 ( .A0(n112), .A1(n2), .A2(n4), .B0(n115), .B1(n113), .Y(n80) );
  NOR2BXL U5 ( .AN(n118), .B(n1), .Y(n122) );
  CLKBUFX3 U6 ( .A(addr[2]), .Y(n4) );
  INVX3 U7 ( .A(addr[6]), .Y(n11) );
  OAI221X4 U8 ( .A0(n88), .A1(n6), .B0(addr[5]), .B1(n87), .C0(n86), .Y(
        dout[2]) );
  OAI221X4 U9 ( .A0(addr[5]), .A1(n127), .B0(n126), .B1(n6), .C0(n125), .Y(
        dout[4]) );
  OA21XL U10 ( .A0(n95), .A1(n115), .B0(n107), .Y(n119) );
  AOI222XL U11 ( .A0(n10), .A1(n1), .B0(n2), .B1(n110), .C0(n12), .C1(n8), .Y(
        n111) );
  AOI2BB2X1 U12 ( .B0(n2), .B1(n12), .A0N(addr[4]), .A1N(n115), .Y(n91) );
  BUFX4 U14 ( .A(addr[3]), .Y(n3) );
  CLKINVX1 U15 ( .A(n112), .Y(n10) );
  CLKINVX1 U16 ( .A(n113), .Y(n7) );
  NAND2BX1 U17 ( .AN(n104), .B(n119), .Y(n84) );
  CLKXOR2X2 U18 ( .A(n72), .B(n8), .Y(n90) );
  NOR2X1 U19 ( .A(n71), .B(n72), .Y(n118) );
  OAI21XL U20 ( .A0(n72), .A1(n114), .B0(n91), .Y(n92) );
  NAND2X1 U21 ( .A(n93), .B(n71), .Y(n107) );
  NAND2X1 U22 ( .A(n8), .B(n72), .Y(n113) );
  OAI211X1 U23 ( .A0(n71), .A1(n114), .B0(n108), .C0(n107), .Y(n89) );
  CLKINVX1 U24 ( .A(n109), .Y(n12) );
  NAND2X1 U25 ( .A(n124), .B(n69), .Y(n108) );
  CLKINVX1 U26 ( .A(n114), .Y(n9) );
  CLKINVX1 U27 ( .A(n115), .Y(n69) );
  CLKINVX1 U28 ( .A(n95), .Y(n5) );
  AO22X1 U29 ( .A0(n90), .A1(n69), .B0(n72), .B1(n123), .Y(n76) );
  OAI31X1 U30 ( .A0(n8), .A1(n3), .A2(n70), .B0(n103), .Y(n105) );
  AOI31XL U31 ( .A0(n70), .A1(n8), .A2(n2), .B0(n102), .Y(n103) );
  AOI211X1 U32 ( .A0(n13), .A1(n4), .B0(n117), .C0(n116), .Y(n126) );
  CLKINVX1 U33 ( .A(n108), .Y(n13) );
  AOI211X1 U34 ( .A0(n115), .A1(n114), .B0(n113), .C0(n2), .Y(n116) );
  OAI22X1 U35 ( .A0(n120), .A1(n112), .B0(n111), .B1(n72), .Y(n117) );
  AOI211X1 U36 ( .A0(n12), .A1(n118), .B0(n81), .C0(n80), .Y(n88) );
  OAI22X1 U37 ( .A0(n91), .A1(n8), .B0(n3), .B1(n106), .Y(n81) );
  CLKINVX3 U38 ( .A(addr[5]), .Y(n6) );
  NAND2X1 U39 ( .A(n3), .B(n6), .Y(n95) );
  NAND2X1 U40 ( .A(n9), .B(n1), .Y(n106) );
  XOR2X1 U41 ( .A(n82), .B(n2), .Y(n83) );
  NAND2X1 U43 ( .A(n1), .B(n3), .Y(n82) );
  OAI22XL U45 ( .A0(n3), .A1(n70), .B0(n72), .B1(n112), .Y(n94) );
  AOI211XL U46 ( .A0(n98), .A1(n72), .B0(n97), .C0(n104), .Y(n99) );
  OAI22XL U47 ( .A0(n96), .A1(n71), .B0(n95), .B1(n109), .Y(n97) );
  OAI22XL U52 ( .A0(n11), .A1(n6), .B0(n2), .B1(addr[1]), .Y(n98) );
  AOI221XL U53 ( .A0(n5), .A1(addr[6]), .B0(addr[5]), .B1(n94), .C0(n93), .Y(
        n96) );
  OAI21XL U54 ( .A0(addr[1]), .A1(n120), .B0(n119), .Y(n121) );
  AOI221XL U58 ( .A0(n10), .A1(n118), .B0(n93), .B1(n6), .C0(n75), .Y(n78) );
  OAI31X1 U60 ( .A0(n6), .A1(n2), .A2(n74), .B0(n73), .Y(n75) );
  OA21XL U61 ( .A0(n3), .A1(n11), .B0(n109), .Y(n74) );
  OAI21XL U62 ( .A0(n124), .A1(n85), .B0(n9), .Y(n73) );
  OAI21XL U63 ( .A0(n1), .A1(n70), .B0(n109), .Y(n110) );
  INVX4 U64 ( .A(n4), .Y(n8) );
  AOI222XL U65 ( .A0(n124), .A1(n123), .B0(n122), .B1(addr[6]), .C0(n1), .C1(
        n121), .Y(n125) );
  NOR4BBX1 U66 ( .AN(n107), .BN(n106), .C(n105), .D(n104), .Y(n127) );
  AOI222XL U67 ( .A0(n10), .A1(n90), .B0(n89), .B1(n8), .C0(n123), .C1(n71), 
        .Y(n101) );
  AOI2BB2XL U68 ( .B0(addr[5]), .B1(n92), .A0N(n120), .A1N(addr[1]), .Y(n100)
         );
  AOI32X1 U69 ( .A0(n4), .A1(n85), .A2(n10), .B0(n84), .B1(n8), .Y(n86) );
  AOI222XL U70 ( .A0(n124), .A1(n70), .B0(n83), .B1(addr[1]), .C0(n7), .C1(n11), .Y(n87) );
  OAI221X1 U71 ( .A0(n79), .A1(n6), .B0(n4), .B1(n78), .C0(n77), .Y(dout[1])
         );
  AOI32XL U72 ( .A0(addr[6]), .A1(n85), .A2(n1), .B0(n76), .B1(n6), .Y(n77) );
  AOI221X1 U73 ( .A0(n10), .A1(n90), .B0(n4), .B1(n93), .C0(n102), .Y(n79) );
  CLKINVX3 U74 ( .A(addr[1]), .Y(n70) );
  CLKINVX3 U75 ( .A(n2), .Y(n71) );
  CLKINVX3 U76 ( .A(n3), .Y(n72) );
endmodule


module sbox2_9 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147;

  NAND2X2 U55 ( .A(n2), .B(n82), .Y(n136) );
  NAND2X2 U57 ( .A(addr[2]), .B(n5), .Y(n104) );
  NAND2X2 U60 ( .A(addr[5]), .B(addr[2]), .Y(n132) );
  NOR2X2 U61 ( .A(n10), .B(n8), .Y(n101) );
  NAND2X2 U62 ( .A(n83), .B(n9), .Y(n146) );
  NAND2X2 U63 ( .A(n3), .B(n13), .Y(n124) );
  NAND2X2 U64 ( .A(addr[6]), .B(n83), .Y(n122) );
  NAND2X2 U67 ( .A(n3), .B(n2), .Y(n133) );
  AOI222XL U1 ( .A0(n14), .A1(n7), .B0(n88), .B1(n13), .C0(n140), .C1(n8), .Y(
        n89) );
  CLKINVX1 U2 ( .A(n121), .Y(n10) );
  CLKINVX1 U3 ( .A(addr[5]), .Y(n1) );
  INVX3 U4 ( .A(addr[5]), .Y(n5) );
  OAI211X4 U5 ( .A0(n147), .A1(n146), .B0(n145), .C0(n144), .Y(dout[4]) );
  NAND3XL U6 ( .A(n98), .B(n97), .C(n96), .Y(dout[1]) );
  NOR2X1 U7 ( .A(n104), .B(n2), .Y(n141) );
  NOR2X1 U8 ( .A(n124), .B(n2), .Y(n140) );
  CLKBUFX4 U9 ( .A(addr[4]), .Y(n2) );
  NAND2X1 U10 ( .A(addr[1]), .B(addr[6]), .Y(n121) );
  CLKINVX2 U11 ( .A(addr[1]), .Y(n83) );
  OAI221X1 U12 ( .A0(addr[1]), .A1(n136), .B0(n133), .B1(n83), .C0(n87), .Y(
        n95) );
  NAND2X4 U13 ( .A(addr[1]), .B(n9), .Y(n114) );
  INVX3 U14 ( .A(addr[6]), .Y(n9) );
  NAND2XL U15 ( .A(n102), .B(n82), .Y(n109) );
  AOI211XL U16 ( .A0(n6), .A1(n95), .B0(n94), .C0(n93), .Y(n96) );
  AOI2BB2X1 U17 ( .B0(n5), .B1(n12), .A0N(n104), .A1N(n136), .Y(n117) );
  NOR3BXL U18 ( .AN(n135), .B(n134), .C(n14), .Y(n147) );
  BUFX4 U19 ( .A(addr[3]), .Y(n3) );
  NAND2X1 U20 ( .A(n14), .B(n10), .Y(n113) );
  CLKINVX1 U21 ( .A(n146), .Y(n8) );
  CLKINVX1 U22 ( .A(n115), .Y(n14) );
  CLKINVX1 U23 ( .A(n122), .Y(n11) );
  OAI31X1 U24 ( .A0(n124), .A1(n9), .A2(n5), .B0(n123), .Y(n128) );
  OAI21XL U25 ( .A0(n5), .A1(n83), .B0(n140), .Y(n123) );
  OAI22X1 U26 ( .A0(n122), .A1(n124), .B0(n101), .B1(n132), .Y(n84) );
  INVX1 U27 ( .A(n114), .Y(n7) );
  OAI22X1 U28 ( .A0(n122), .A1(n82), .B0(n15), .B1(n121), .Y(n129) );
  NAND3X1 U29 ( .A(n15), .B(n5), .C(n83), .Y(n111) );
  NAND2X1 U30 ( .A(n82), .B(n15), .Y(n115) );
  OAI21XL U31 ( .A0(n13), .A1(n133), .B0(n135), .Y(n85) );
  OAI22XL U32 ( .A0(n117), .A1(n146), .B0(n116), .B1(n132), .Y(n118) );
  AOI222XL U33 ( .A0(n7), .A1(n115), .B0(n16), .B1(n9), .C0(n14), .C1(n8), .Y(
        n116) );
  CLKINVX1 U34 ( .A(n104), .Y(n4) );
  OAI2BB2XL U35 ( .B0(n114), .B1(n135), .A0N(n126), .A1N(n16), .Y(n106) );
  OAI21XL U36 ( .A0(n112), .A1(n114), .B0(n111), .Y(n120) );
  OAI21XL U37 ( .A0(n133), .A1(n114), .B0(n113), .Y(n119) );
  CLKINVX1 U38 ( .A(n124), .Y(n12) );
  CLKINVX1 U39 ( .A(n136), .Y(n81) );
  CLKINVX1 U40 ( .A(n133), .Y(n16) );
  CLKINVX1 U41 ( .A(n132), .Y(n6) );
  AOI2BB1X1 U42 ( .A0N(n126), .A1N(n125), .B0(n136), .Y(n127) );
  OAI22XL U43 ( .A0(n104), .A1(n114), .B0(n101), .B1(n132), .Y(n102) );
  AO21XL U44 ( .A0(n13), .A1(n81), .B0(n141), .Y(n86) );
  AO21X1 U45 ( .A0(n82), .A1(n4), .B0(n140), .Y(n142) );
  NAND3X1 U46 ( .A(n13), .B(n15), .C(addr[5]), .Y(n135) );
  OAI22X1 U47 ( .A0(addr[5]), .A1(n121), .B0(n122), .B1(n5), .Y(n126) );
  AOI2BB1X1 U48 ( .A0N(n3), .A1N(n1), .B0(n81), .Y(n112) );
  NOR3X1 U49 ( .A(addr[1]), .B(addr[2]), .C(n5), .Y(n125) );
  AOI2BB1XL U50 ( .A0N(n92), .A1N(n91), .B0(addr[5]), .Y(n93) );
  OAI22XL U51 ( .A0(n117), .A1(n114), .B0(n89), .B1(n1), .Y(n94) );
  OAI31XL U52 ( .A0(n114), .A1(n2), .A2(n82), .B0(n90), .Y(n91) );
  OAI21XL U53 ( .A0(n16), .A1(n12), .B0(n11), .Y(n90) );
  NAND2X1 U54 ( .A(n7), .B(n2), .Y(n137) );
  OAI31XL U56 ( .A0(n101), .A1(n3), .A2(addr[2]), .B0(n113), .Y(n92) );
  OAI211X1 U58 ( .A0(n139), .A1(n5), .B0(n138), .C0(n137), .Y(n143) );
  NAND3X1 U59 ( .A(n15), .B(n5), .C(addr[6]), .Y(n138) );
  AOI2BB2X1 U65 ( .B0(n11), .B1(n82), .A0N(n83), .A1N(n136), .Y(n139) );
  OAI22XL U66 ( .A0(addr[5]), .A1(n133), .B0(n3), .B1(n132), .Y(n134) );
  OAI2BB2XL U68 ( .B0(n112), .B1(n122), .A0N(n1), .A1N(n99), .Y(n100) );
  OAI211X1 U69 ( .A0(n146), .A1(n2), .B0(n137), .C0(n113), .Y(n99) );
  NAND3X1 U70 ( .A(n11), .B(n15), .C(n3), .Y(n87) );
  AOI2BB2XL U71 ( .B0(n3), .B1(n105), .A0N(n137), .A1N(n132), .Y(n108) );
  OAI211XL U72 ( .A0(n104), .A1(n146), .B0(n103), .C0(n111), .Y(n105) );
  NAND3XL U73 ( .A(addr[5]), .B(n15), .C(n10), .Y(n103) );
  OAI22XL U74 ( .A0(n3), .A1(n114), .B0(n9), .B1(n115), .Y(n88) );
  NAND4X1 U75 ( .A(n110), .B(n109), .C(n108), .D(n107), .Y(dout[2]) );
  AOI32XL U76 ( .A0(addr[1]), .A1(addr[2]), .A2(n81), .B0(n100), .B1(n13), .Y(
        n110) );
  AOI221XL U77 ( .A0(n125), .A1(addr[4]), .B0(n141), .B1(n11), .C0(n106), .Y(
        n107) );
  AOI33XL U78 ( .A0(n11), .A1(n4), .A2(n2), .B0(n6), .B1(n146), .B2(n3), .Y(
        n145) );
  AOI222XL U79 ( .A0(n143), .A1(n13), .B0(n10), .B1(n142), .C0(n7), .C1(n141), 
        .Y(n144) );
  AOI32XL U80 ( .A0(n4), .A1(n83), .A2(n14), .B0(n8), .B1(n86), .Y(n97) );
  AOI22X1 U81 ( .A0(n10), .A1(n85), .B0(n2), .B1(n84), .Y(n98) );
  NAND2X1 U82 ( .A(n131), .B(n130), .Y(dout[3]) );
  AOI221XL U83 ( .A0(n120), .A1(n13), .B0(addr[2]), .B1(n119), .C0(n118), .Y(
        n131) );
  AOI211X1 U84 ( .A0(n4), .A1(n129), .B0(n128), .C0(n127), .Y(n130) );
  CLKINVX3 U85 ( .A(addr[2]), .Y(n13) );
  CLKINVX3 U86 ( .A(n2), .Y(n15) );
  CLKINVX3 U87 ( .A(n3), .Y(n82) );
endmodule


module sbox3_9 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134;

  NOR2X2 U35 ( .A(n76), .B(addr[3]), .Y(n109) );
  NOR2X2 U50 ( .A(addr[1]), .B(addr[6]), .Y(n108) );
  NOR2X2 U52 ( .A(n78), .B(n3), .Y(n88) );
  NOR2X2 U56 ( .A(n78), .B(n16), .Y(n95) );
  NOR2X1 U1 ( .A(n76), .B(n78), .Y(n107) );
  OAI221X1 U2 ( .A0(n125), .A1(n76), .B0(n4), .B1(addr[1]), .C0(n14), .Y(n105)
         );
  INVXL U3 ( .A(n2), .Y(n1) );
  NOR2X1 U4 ( .A(n10), .B(n4), .Y(n92) );
  NOR2X1 U5 ( .A(n77), .B(n4), .Y(n122) );
  NOR2X1 U6 ( .A(n14), .B(n4), .Y(n96) );
  CLKBUFX3 U7 ( .A(addr[2]), .Y(n4) );
  INVX1 U8 ( .A(addr[2]), .Y(n2) );
  NOR2X1 U9 ( .A(n4), .B(n3), .Y(n111) );
  BUFX4 U10 ( .A(addr[4]), .Y(n3) );
  OAI33X1 U11 ( .A0(n77), .A1(n126), .A2(n16), .B0(n76), .B1(n95), .B2(n120), 
        .Y(n80) );
  INVX3 U12 ( .A(n4), .Y(n16) );
  OAI221X1 U13 ( .A0(addr[5]), .A1(n91), .B0(n90), .B1(n19), .C0(n89), .Y(
        dout[1]) );
  NOR2X4 U14 ( .A(n11), .B(n79), .Y(n125) );
  NOR2X4 U15 ( .A(addr[3]), .B(n3), .Y(n131) );
  NOR2X4 U16 ( .A(n79), .B(addr[6]), .Y(n126) );
  INVX3 U17 ( .A(addr[1]), .Y(n79) );
  NAND2XL U18 ( .A(n95), .B(n125), .Y(n133) );
  OAI211XL U19 ( .A0(n3), .A1(n9), .B0(n129), .C0(n128), .Y(n130) );
  NAND4XL U20 ( .A(n115), .B(n114), .C(n113), .D(n112), .Y(n116) );
  CLKINVX1 U21 ( .A(n133), .Y(n7) );
  INVX1 U22 ( .A(n125), .Y(n5) );
  CLKINVX1 U23 ( .A(n107), .Y(n20) );
  NAND2X1 U24 ( .A(n10), .B(n12), .Y(n123) );
  CLKINVX1 U25 ( .A(n87), .Y(n12) );
  CLKINVX1 U26 ( .A(n121), .Y(n15) );
  CLKINVX1 U27 ( .A(n120), .Y(n6) );
  CLKINVX1 U28 ( .A(n115), .Y(n8) );
  CLKINVX1 U29 ( .A(n108), .Y(n14) );
  NOR2X1 U30 ( .A(n10), .B(n16), .Y(n104) );
  NOR2X1 U31 ( .A(n5), .B(n16), .Y(n110) );
  INVX1 U32 ( .A(n126), .Y(n13) );
  AOI21X1 U33 ( .A0(n78), .A1(n16), .B0(n95), .Y(n121) );
  OAI21XL U34 ( .A0(n111), .A1(n131), .B0(n125), .Y(n83) );
  CLKINVX1 U36 ( .A(n82), .Y(n10) );
  NOR2X1 U37 ( .A(n13), .B(n76), .Y(n87) );
  NOR2X1 U38 ( .A(n125), .B(n108), .Y(n120) );
  OAI21XL U39 ( .A0(n110), .A1(n92), .B0(n131), .Y(n101) );
  NAND2X1 U40 ( .A(n104), .B(n88), .Y(n115) );
  CLKINVX1 U41 ( .A(n88), .Y(n77) );
  CLKINVX1 U42 ( .A(n92), .Y(n9) );
  CLKINVX1 U43 ( .A(n111), .Y(n17) );
  CLKINVX1 U44 ( .A(n122), .Y(n18) );
  OR2X1 U45 ( .A(n104), .B(n96), .Y(n127) );
  OAI221X1 U46 ( .A0(n13), .A1(n17), .B0(n16), .B1(n12), .C0(n94), .Y(n99) );
  AOI221XL U47 ( .A0(n96), .A1(n3), .B0(n93), .B1(n76), .C0(n7), .Y(n94) );
  OAI21XL U48 ( .A0(n16), .A1(n14), .B0(n9), .Y(n93) );
  XNOR2X1 U49 ( .A(addr[5]), .B(addr[3]), .Y(n103) );
  CLKINVX1 U51 ( .A(addr[5]), .Y(n19) );
  OAI221X1 U53 ( .A0(n14), .A1(n17), .B0(n5), .B1(n77), .C0(n106), .Y(n117) );
  AOI221XL U54 ( .A0(addr[3]), .A1(n105), .B0(n104), .B1(n131), .C0(n7), .Y(
        n106) );
  CLKINVX1 U55 ( .A(addr[6]), .Y(n11) );
  NAND3X1 U57 ( .A(n4), .B(n79), .C(n109), .Y(n114) );
  NOR2X1 U58 ( .A(n11), .B(addr[1]), .Y(n82) );
  AOI32XL U59 ( .A0(n16), .A1(n78), .A2(n125), .B0(n124), .B1(n11), .Y(n129)
         );
  AOI22XL U60 ( .A0(n3), .A1(n127), .B0(n126), .B1(n131), .Y(n128) );
  OAI22XL U61 ( .A0(n3), .A1(n2), .B0(n4), .B1(n20), .Y(n124) );
  AOI222XL U62 ( .A0(n111), .A1(n126), .B0(n110), .B1(n78), .C0(n109), .C1(
        n108), .Y(n112) );
  OAI211XL U63 ( .A0(n107), .A1(n131), .B0(n2), .C0(addr[6]), .Y(n113) );
  OAI21XL U64 ( .A0(n1), .A1(addr[1]), .B0(n13), .Y(n81) );
  AOI221XL U65 ( .A0(n87), .A1(n78), .B0(n88), .B1(n126), .C0(n86), .Y(n90) );
  OAI211X1 U66 ( .A0(n85), .A1(n16), .B0(n84), .C0(n83), .Y(n86) );
  AOI222XL U67 ( .A0(n82), .A1(n78), .B0(n108), .B1(n107), .C0(n131), .C1(n79), 
        .Y(n85) );
  OAI21XL U68 ( .A0(n92), .A1(n7), .B0(addr[4]), .Y(n84) );
  AOI221XL U69 ( .A0(n126), .A1(n15), .B0(addr[3]), .B1(n127), .C0(n97), .Y(
        n98) );
  OAI22X1 U70 ( .A0(n5), .A1(n18), .B0(n20), .B1(n10), .Y(n97) );
  OAI211X1 U71 ( .A0(n14), .A1(n18), .B0(n119), .C0(n118), .Y(dout[3]) );
  AOI32XL U72 ( .A0(n126), .A1(n4), .A2(n103), .B0(n109), .B1(n110), .Y(n119)
         );
  AOI22XL U73 ( .A0(n117), .A1(n19), .B0(addr[5]), .B1(n116), .Y(n118) );
  AOI221XL U74 ( .A0(n122), .A1(n126), .B0(n96), .B1(n109), .C0(n8), .Y(n89)
         );
  AOI221XL U75 ( .A0(n131), .A1(n81), .B0(n95), .B1(n123), .C0(n80), .Y(n91)
         );
  NAND4X1 U76 ( .A(n102), .B(n114), .C(n101), .D(n100), .Y(dout[2]) );
  NAND3XL U77 ( .A(n3), .B(n125), .C(n103), .Y(n102) );
  AOI2BB2XL U78 ( .B0(addr[5]), .B1(n99), .A0N(addr[5]), .A1N(n98), .Y(n100)
         );
  OAI221X1 U79 ( .A0(n134), .A1(n19), .B0(n3), .B1(n133), .C0(n132), .Y(
        dout[4]) );
  AOI32XL U80 ( .A0(n131), .A1(n11), .A2(n1), .B0(n130), .B1(n19), .Y(n132) );
  AOI222XL U81 ( .A0(n15), .A1(n123), .B0(n122), .B1(addr[1]), .C0(n121), .C1(
        n6), .Y(n134) );
  CLKINVX3 U82 ( .A(n3), .Y(n76) );
  CLKINVX3 U83 ( .A(addr[3]), .Y(n78) );
endmodule


module sbox4_9 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126;

  OAI32X4 U12 ( .A0(n12), .A1(n2), .A2(addr[2]), .B0(n71), .B1(n108), .Y(n123)
         );
  OAI222X4 U20 ( .A0(addr[2]), .A1(n92), .B0(n106), .B1(n91), .C0(n90), .C1(
        n16), .Y(dout[2]) );
  OAI222X4 U33 ( .A0(addr[4]), .A1(n106), .B0(n72), .B1(n108), .C0(n2), .C1(
        n118), .Y(n83) );
  NAND2X2 U34 ( .A(addr[4]), .B(n2), .Y(n108) );
  NOR2X2 U43 ( .A(n14), .B(addr[4]), .Y(n113) );
  NOR2X2 U45 ( .A(n71), .B(n2), .Y(n111) );
  NAND2X2 U51 ( .A(n72), .B(n8), .Y(n118) );
  NOR2X2 U52 ( .A(n13), .B(addr[5]), .Y(n97) );
  NAND2X2 U53 ( .A(addr[6]), .B(addr[1]), .Y(n85) );
  NAND2X2 U54 ( .A(addr[1]), .B(n8), .Y(n116) );
  NOR2X2 U55 ( .A(n115), .B(n71), .Y(n121) );
  NAND2X2 U56 ( .A(n14), .B(n13), .Y(n115) );
  NAND2X2 U57 ( .A(addr[5]), .B(n13), .Y(n96) );
  NAND2X2 U58 ( .A(addr[6]), .B(n72), .Y(n106) );
  OAI222X1 U1 ( .A0(n12), .A1(n85), .B0(n97), .B1(n116), .C0(n13), .C1(n118), 
        .Y(n73) );
  CLKINVX1 U2 ( .A(n116), .Y(n7) );
  CLKINVX1 U3 ( .A(n14), .Y(n1) );
  CLKBUFX3 U4 ( .A(addr[3]), .Y(n2) );
  OAI31X4 U5 ( .A0(n118), .A1(n71), .A2(n13), .B0(n117), .Y(n119) );
  OAI221X1 U6 ( .A0(addr[2]), .A1(n80), .B0(n118), .B1(n105), .C0(n79), .Y(
        dout[1]) );
  AOI222XL U7 ( .A0(n13), .A1(n8), .B0(n113), .B1(n72), .C0(addr[1]), .C1(n14), 
        .Y(n114) );
  OAI222X1 U8 ( .A0(addr[1]), .A1(n84), .B0(n85), .B1(n74), .C0(n14), .C1(n107), .Y(n75) );
  INVX4 U9 ( .A(addr[5]), .Y(n71) );
  OAI31X1 U10 ( .A0(n108), .A1(addr[5]), .A2(n9), .B0(n107), .Y(n109) );
  NAND2XL U11 ( .A(n1), .B(addr[5]), .Y(n84) );
  AOI211XL U13 ( .A0(n83), .A1(n71), .B0(n82), .C0(n4), .Y(n92) );
  NAND2XL U14 ( .A(n13), .B(n71), .Y(n74) );
  CLKINVX1 U15 ( .A(n118), .Y(n3) );
  CLKINVX1 U16 ( .A(n115), .Y(n11) );
  CLKINVX1 U17 ( .A(n112), .Y(n6) );
  OAI21X1 U18 ( .A0(n7), .A1(n9), .B0(n16), .Y(n112) );
  AOI22X1 U19 ( .A0(n10), .A1(n111), .B0(n9), .B1(n113), .Y(n93) );
  OAI211X1 U21 ( .A0(n72), .A1(n115), .B0(n93), .C0(n5), .Y(n94) );
  CLKINVX1 U22 ( .A(n85), .Y(n10) );
  NAND2X1 U23 ( .A(n97), .B(n14), .Y(n105) );
  NAND2X1 U24 ( .A(n113), .B(n3), .Y(n98) );
  NAND2X1 U25 ( .A(n7), .B(n97), .Y(n107) );
  NAND2X1 U26 ( .A(n118), .B(n85), .Y(n110) );
  OAI21XL U27 ( .A0(n11), .A1(n71), .B0(n108), .Y(n95) );
  CLKINVX1 U28 ( .A(n84), .Y(n15) );
  CLKINVX1 U29 ( .A(addr[2]), .Y(n16) );
  OAI31X1 U30 ( .A0(n13), .A1(addr[6]), .A2(n71), .B0(n87), .Y(n88) );
  OAI21XL U31 ( .A0(n113), .A1(n12), .B0(n10), .Y(n87) );
  OAI211X1 U32 ( .A0(n76), .A1(n13), .B0(n98), .C0(n5), .Y(n77) );
  AOI222XL U35 ( .A0(addr[5]), .A1(addr[6]), .B0(n111), .B1(addr[1]), .C0(n9), 
        .C1(n2), .Y(n76) );
  NAND3XL U36 ( .A(n10), .B(n14), .C(addr[4]), .Y(n117) );
  OAI22XL U37 ( .A0(n116), .A1(n115), .B0(n1), .B1(n112), .Y(n78) );
  CLKINVX3 U38 ( .A(addr[4]), .Y(n13) );
  OAI2BB2XL U39 ( .B0(n115), .B1(n106), .A0N(n71), .A1N(n86), .Y(n89) );
  OAI221XL U40 ( .A0(n116), .A1(addr[4]), .B0(n108), .B1(addr[1]), .C0(n117), 
        .Y(n86) );
  CLKINVX1 U41 ( .A(addr[6]), .Y(n8) );
  CLKINVX1 U42 ( .A(n81), .Y(n4) );
  OAI21XL U44 ( .A0(n96), .A1(n118), .B0(n93), .Y(n82) );
  NAND3X1 U46 ( .A(n101), .B(n100), .C(n99), .Y(n102) );
  AOI32X1 U47 ( .A0(n96), .A1(n14), .A2(n7), .B0(n10), .B1(n95), .Y(n101) );
  AOI2BB2XL U48 ( .B0(n72), .B1(n121), .A0N(n98), .A1N(addr[5]), .Y(n99) );
  OAI21XL U49 ( .A0(n97), .A1(n12), .B0(n9), .Y(n100) );
  AOI2BB2XL U50 ( .B0(n9), .B1(n123), .A0N(n122), .A1N(n16), .Y(n124) );
  AOI211XL U59 ( .A0(n9), .A1(n121), .B0(n120), .C0(n119), .Y(n122) );
  OAI22XL U60 ( .A0(n116), .A1(n115), .B0(addr[5]), .B1(n114), .Y(n120) );
  CLKINVX1 U61 ( .A(n75), .Y(n5) );
  AOI32XL U62 ( .A0(n7), .A1(n96), .A2(n1), .B0(addr[1]), .B1(n121), .Y(n81)
         );
  AOI222XL U63 ( .A0(n9), .A1(n12), .B0(n121), .B1(n116), .C0(n2), .C1(n73), 
        .Y(n80) );
  AOI22XL U64 ( .A0(n78), .A1(n71), .B0(addr[2]), .B1(n77), .Y(n79) );
  NAND2XL U65 ( .A(n111), .B(addr[4]), .Y(n91) );
  AOI211X1 U66 ( .A0(n15), .A1(n110), .B0(n89), .C0(n88), .Y(n90) );
  OAI211X1 U67 ( .A0(n106), .A1(n105), .B0(n104), .C0(n103), .Y(dout[3]) );
  AOI32X1 U68 ( .A0(n2), .A1(n12), .A2(n7), .B0(n94), .B1(n16), .Y(n104) );
  AOI22XL U69 ( .A0(addr[2]), .A1(n102), .B0(n3), .B1(n123), .Y(n103) );
  OAI211X1 U70 ( .A0(addr[2]), .A1(n126), .B0(n125), .C0(n124), .Y(dout[4]) );
  AOI32X1 U71 ( .A0(n10), .A1(n12), .A2(n2), .B0(n6), .B1(n15), .Y(n125) );
  AOI221XL U72 ( .A0(n3), .A1(n111), .B0(n11), .B1(n110), .C0(n109), .Y(n126)
         );
  CLKINVX3 U73 ( .A(n106), .Y(n9) );
  CLKINVX3 U74 ( .A(n96), .Y(n12) );
  CLKINVX3 U75 ( .A(n2), .Y(n14) );
  CLKINVX3 U76 ( .A(addr[1]), .Y(n72) );
endmodule


module sbox5_9 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121;

  OAI222X4 U18 ( .A0(addr[3]), .A1(n106), .B0(n13), .B1(n90), .C0(n16), .C1(n8), .Y(n93) );
  OAI22X2 U40 ( .A0(addr[5]), .A1(n106), .B0(n14), .B1(n114), .Y(n116) );
  NOR2X2 U41 ( .A(n3), .B(addr[3]), .Y(n102) );
  NAND2X2 U45 ( .A(addr[6]), .B(n8), .Y(n114) );
  NAND2X2 U50 ( .A(n8), .B(n13), .Y(n110) );
  NAND2X2 U52 ( .A(addr[1]), .B(n13), .Y(n113) );
  NAND2X2 U54 ( .A(addr[1]), .B(addr[6]), .Y(n106) );
  NAND2X2 U55 ( .A(addr[3]), .B(n16), .Y(n121) );
  OAI31X1 U1 ( .A0(n70), .A1(addr[5]), .A2(addr[1]), .B0(n81), .Y(n73) );
  CLKINVX1 U2 ( .A(addr[5]), .Y(n1) );
  AOI221XL U3 ( .A0(n93), .A1(n1), .B0(n9), .B1(n68), .C0(n92), .Y(n105) );
  INVX3 U4 ( .A(addr[5]), .Y(n14) );
  OAI221X4 U5 ( .A0(n111), .A1(n110), .B0(n121), .B1(n114), .C0(n109), .Y(n112) );
  OAI221X4 U6 ( .A0(n16), .A1(n114), .B0(n14), .B1(n113), .C0(n120), .Y(n115)
         );
  OAI221X4 U7 ( .A0(n107), .A1(n121), .B0(n111), .B1(n113), .C0(n85), .Y(n86)
         );
  OAI32X1 U8 ( .A0(n114), .A1(addr[5]), .A2(n3), .B0(n15), .B1(n107), .Y(n79)
         );
  AOI32XL U9 ( .A0(n68), .A1(n98), .A2(n11), .B0(n2), .B1(n73), .Y(n77) );
  CLKBUFX3 U10 ( .A(addr[4]), .Y(n2) );
  CLKINVX1 U11 ( .A(n81), .Y(n4) );
  NAND2X1 U12 ( .A(n5), .B(n68), .Y(n81) );
  CLKINVX1 U13 ( .A(n110), .Y(n7) );
  CLKXOR2X2 U14 ( .A(n70), .B(n14), .Y(n94) );
  AOI2BB1X1 U15 ( .A0N(n16), .A1N(n1), .B0(n68), .Y(n111) );
  NOR2X1 U16 ( .A(n121), .B(n14), .Y(n91) );
  NOR2BX1 U17 ( .AN(n116), .B(n90), .Y(n83) );
  NAND2X1 U19 ( .A(n7), .B(n14), .Y(n120) );
  CLKINVX1 U20 ( .A(n113), .Y(n11) );
  NAND2X1 U21 ( .A(n11), .B(n14), .Y(n107) );
  CLKINVX1 U22 ( .A(n121), .Y(n15) );
  OAI31X1 U23 ( .A0(n12), .A1(n68), .A2(n113), .B0(n99), .Y(n72) );
  CLKINVX1 U24 ( .A(n106), .Y(n9) );
  OAI2BB2XL U25 ( .B0(n1), .B1(n113), .A0N(n98), .A1N(n5), .Y(n101) );
  CLKINVX1 U26 ( .A(n114), .Y(n5) );
  CLKINVX1 U27 ( .A(n90), .Y(n69) );
  CLKINVX1 U28 ( .A(addr[1]), .Y(n8) );
  CLKINVX1 U29 ( .A(addr[3]), .Y(n70) );
  CLKINVX1 U30 ( .A(addr[6]), .Y(n13) );
  AOI211X1 U31 ( .A0(n91), .A1(addr[1]), .B0(n80), .C0(n79), .Y(n89) );
  OAI2BB2XL U32 ( .B0(n111), .B1(n106), .A0N(n94), .A1N(n7), .Y(n80) );
  AOI211X1 U33 ( .A0(n102), .A1(n84), .B0(n83), .C0(n82), .Y(n85) );
  OAI21XL U34 ( .A0(n13), .A1(n1), .B0(n106), .Y(n84) );
  NOR3XL U35 ( .A(n94), .B(n3), .C(n110), .Y(n82) );
  AOI222XL U36 ( .A0(n9), .A1(n69), .B0(addr[5]), .B1(n108), .C0(n10), .C1(n16), .Y(n109) );
  CLKINVX1 U37 ( .A(n107), .Y(n10) );
  OAI21XL U38 ( .A0(addr[6]), .A1(addr[3]), .B0(n106), .Y(n108) );
  NAND2X1 U39 ( .A(addr[3]), .B(n3), .Y(n90) );
  NAND2X1 U42 ( .A(n2), .B(addr[5]), .Y(n98) );
  NAND2X1 U43 ( .A(n3), .B(n70), .Y(n97) );
  OAI21XL U44 ( .A0(addr[1]), .A1(n97), .B0(n96), .Y(n103) );
  AOI33XL U46 ( .A0(n3), .A1(n95), .A2(addr[5]), .B0(n94), .B1(n16), .B2(
        addr[1]), .Y(n96) );
  OAI21XL U47 ( .A0(n8), .A1(n70), .B0(n114), .Y(n95) );
  OAI21XL U48 ( .A0(addr[6]), .A1(n121), .B0(n99), .Y(n100) );
  NAND2X1 U49 ( .A(n71), .B(n7), .Y(n99) );
  XOR2X1 U51 ( .A(n12), .B(n3), .Y(n71) );
  AOI2BB2XL U53 ( .B0(n102), .B1(n116), .A0N(n2), .A1N(n75), .Y(n76) );
  AOI211X1 U56 ( .A0(n6), .A1(n3), .B0(n74), .C0(n83), .Y(n75) );
  AO22XL U57 ( .A0(n11), .A1(n15), .B0(addr[6]), .B1(n102), .Y(n74) );
  CLKINVX1 U58 ( .A(n120), .Y(n6) );
  CLKINVX1 U59 ( .A(n2), .Y(n12) );
  AO22XL U60 ( .A0(n11), .A1(n69), .B0(addr[6]), .B1(n91), .Y(n92) );
  AOI222XL U61 ( .A0(n116), .A1(n16), .B0(addr[3]), .B1(n115), .C0(n11), .C1(
        n68), .Y(n117) );
  OAI221X1 U62 ( .A0(n2), .A1(n105), .B0(n110), .B1(n121), .C0(n104), .Y(
        dout[3]) );
  AOI222XL U63 ( .A0(n2), .A1(n103), .B0(n102), .B1(n101), .C0(n100), .C1(n1), 
        .Y(n104) );
  OAI211X1 U64 ( .A0(n2), .A1(n89), .B0(n88), .C0(n87), .Y(dout[2]) );
  AOI33XL U65 ( .A0(n15), .A1(n98), .A2(n5), .B0(n3), .B1(n94), .B2(n7), .Y(
        n88) );
  AOI222XL U66 ( .A0(n4), .A1(n14), .B0(n2), .B1(n86), .C0(n91), .C1(n9), .Y(
        n87) );
  OAI211X1 U67 ( .A0(n78), .A1(n14), .B0(n77), .C0(n76), .Y(dout[1]) );
  AOI221XL U68 ( .A0(n15), .A1(addr[1]), .B0(n9), .B1(n68), .C0(n72), .Y(n78)
         );
  OAI211X1 U69 ( .A0(n121), .A1(n120), .B0(n119), .C0(n118), .Y(dout[4]) );
  AOI32XL U70 ( .A0(n68), .A1(n114), .A2(addr[5]), .B0(n2), .B1(n112), .Y(n119) );
  AOI2BB2X1 U71 ( .B0(n4), .B1(n14), .A0N(n2), .A1N(n117), .Y(n118) );
  BUFX4 U72 ( .A(addr[2]), .Y(n3) );
  CLKINVX3 U73 ( .A(n3), .Y(n16) );
  CLKINVX3 U74 ( .A(n97), .Y(n68) );
endmodule


module sbox6_9 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147;

  NAND2X2 U39 ( .A(n138), .B(addr[3]), .Y(n147) );
  NOR2X2 U47 ( .A(n15), .B(n10), .Y(n138) );
  NOR2X2 U50 ( .A(n85), .B(n4), .Y(n119) );
  NOR2X2 U58 ( .A(n83), .B(n85), .Y(n125) );
  NAND2X2 U61 ( .A(n97), .B(n103), .Y(n112) );
  NOR2X2 U62 ( .A(n17), .B(addr[1]), .Y(n103) );
  NOR2X2 U63 ( .A(n83), .B(addr[3]), .Y(n97) );
  NAND2X2 U64 ( .A(n117), .B(n131), .Y(n140) );
  NOR2X2 U65 ( .A(n5), .B(addr[3]), .Y(n131) );
  NOR2X2 U66 ( .A(n11), .B(addr[6]), .Y(n117) );
  NOR2X1 U1 ( .A(n15), .B(addr[3]), .Y(n102) );
  AOI211X1 U2 ( .A0(n18), .A1(n85), .B0(n131), .C0(n143), .Y(n121) );
  CLKINVX1 U3 ( .A(n15), .Y(n1) );
  OAI222X1 U4 ( .A0(n91), .A1(n18), .B0(n5), .B1(n82), .C0(addr[5]), .C1(n84), 
        .Y(n92) );
  BUFX4 U5 ( .A(addr[2]), .Y(n5) );
  CLKINVX1 U6 ( .A(n83), .Y(n2) );
  INVX4 U7 ( .A(n4), .Y(n83) );
  CLKBUFX3 U8 ( .A(addr[4]), .Y(n4) );
  OAI221X1 U9 ( .A0(n17), .A1(n81), .B0(n85), .B1(n8), .C0(n86), .Y(n90) );
  INVX2 U10 ( .A(n96), .Y(n8) );
  CLKINVX1 U11 ( .A(addr[3]), .Y(n3) );
  INVX3 U12 ( .A(addr[3]), .Y(n85) );
  OAI221X4 U13 ( .A0(n123), .A1(n13), .B0(n10), .B1(n18), .C0(n7), .Y(n124) );
  NOR2X4 U14 ( .A(addr[1]), .B(addr[6]), .Y(n130) );
  NOR2X4 U15 ( .A(n5), .B(addr[5]), .Y(n143) );
  INVX1 U16 ( .A(n130), .Y(n14) );
  CLKINVX1 U17 ( .A(n125), .Y(n81) );
  NAND2X1 U18 ( .A(n14), .B(n8), .Y(n105) );
  INVXL U19 ( .A(n121), .Y(n16) );
  CLKINVX1 U20 ( .A(n138), .Y(n9) );
  CLKINVX1 U21 ( .A(n117), .Y(n10) );
  CLKINVX1 U22 ( .A(n119), .Y(n84) );
  NOR2X1 U23 ( .A(n8), .B(n123), .Y(n144) );
  NOR2X1 U24 ( .A(n11), .B(n17), .Y(n96) );
  CLKINVX1 U25 ( .A(n103), .Y(n13) );
  OAI211X1 U26 ( .A0(n14), .A1(n81), .B0(n104), .C0(n112), .Y(n108) );
  OAI21XL U27 ( .A0(n103), .A1(n117), .B0(n102), .Y(n104) );
  OAI21XL U28 ( .A0(n132), .A1(n17), .B0(n3), .Y(n86) );
  AOI21X1 U29 ( .A0(n83), .A1(n102), .B0(n125), .Y(n91) );
  OAI2BB2XL U30 ( .B0(n143), .B1(n14), .A0N(n143), .A1N(n117), .Y(n118) );
  CLKINVX1 U31 ( .A(n122), .Y(n7) );
  CLKINVX1 U32 ( .A(n126), .Y(n12) );
  CLKINVX1 U33 ( .A(n97), .Y(n82) );
  NAND2BX1 U34 ( .AN(n144), .B(n137), .Y(n107) );
  CLKINVX1 U35 ( .A(addr[1]), .Y(n11) );
  NOR2X1 U36 ( .A(n8), .B(n1), .Y(n122) );
  NOR2X1 U37 ( .A(addr[1]), .B(n2), .Y(n132) );
  OAI22X1 U38 ( .A0(n84), .A1(n10), .B0(n5), .B1(n12), .Y(n88) );
  NAND2X1 U40 ( .A(n1), .B(n18), .Y(n123) );
  NAND4X1 U41 ( .A(n147), .B(n140), .C(n100), .D(n99), .Y(n101) );
  AOI222XL U42 ( .A0(n98), .A1(n15), .B0(n102), .B1(n130), .C0(n97), .C1(n105), 
        .Y(n99) );
  NAND3X1 U43 ( .A(n5), .B(n84), .C(n96), .Y(n100) );
  OAI221X1 U44 ( .A0(n85), .A1(n13), .B0(n84), .B1(n17), .C0(n12), .Y(n98) );
  AOI22X1 U45 ( .A0(n4), .A1(n115), .B0(addr[5]), .B1(n114), .Y(n129) );
  OAI21XL U46 ( .A0(n121), .A1(n14), .B0(n147), .Y(n115) );
  OAI21XL U48 ( .A0(n113), .A1(n15), .B0(n112), .Y(n114) );
  AOI221XL U49 ( .A0(n119), .A1(n11), .B0(n130), .B1(addr[3]), .C0(n111), .Y(
        n113) );
  OAI22XL U51 ( .A0(n10), .A1(n83), .B0(addr[3]), .B1(n8), .Y(n111) );
  OAI22XL U52 ( .A0(n85), .A1(n17), .B0(addr[1]), .B1(n84), .Y(n142) );
  AOI211X1 U53 ( .A0(n4), .A1(n135), .B0(n134), .C0(n133), .Y(n136) );
  OA21XL U54 ( .A0(n3), .A1(n1), .B0(n132), .Y(n133) );
  OAI2BB2XL U55 ( .B0(n2), .B1(n7), .A0N(n131), .A1N(n130), .Y(n134) );
  OAI22X1 U56 ( .A0(n5), .A1(n10), .B0(n15), .B1(n8), .Y(n135) );
  CLKINVX3 U57 ( .A(addr[5]), .Y(n18) );
  AOI2BB2X1 U59 ( .B0(n5), .B1(n130), .A0N(n1), .A1N(n13), .Y(n137) );
  NOR2X1 U60 ( .A(n13), .B(n2), .Y(n126) );
  AOI2BB2XL U67 ( .B0(n143), .B1(n90), .A0N(n89), .A1N(n18), .Y(n94) );
  AOI211X1 U68 ( .A0(n122), .A1(n4), .B0(n88), .C0(n87), .Y(n89) );
  OAI32X1 U69 ( .A0(n13), .A1(n85), .A2(n15), .B0(n9), .B1(n82), .Y(n87) );
  NAND3X1 U70 ( .A(n147), .B(n140), .C(n139), .Y(n141) );
  AOI32X1 U71 ( .A0(n5), .A1(n11), .A2(n4), .B0(n138), .B1(n83), .Y(n139) );
  AO22XL U72 ( .A0(n143), .A1(n2), .B0(n116), .B1(n83), .Y(n120) );
  OAI21XL U73 ( .A0(n1), .A1(n18), .B0(n123), .Y(n116) );
  CLKINVX1 U74 ( .A(n106), .Y(n6) );
  AOI32XL U75 ( .A0(n105), .A1(n83), .A2(n3), .B0(addr[1]), .B1(n125), .Y(n106) );
  OAI211X1 U76 ( .A0(n83), .A1(n140), .B0(n110), .C0(n109), .Y(dout[2]) );
  AOI222XL U77 ( .A0(n108), .A1(n18), .B0(n143), .B1(n6), .C0(n119), .C1(n107), 
        .Y(n109) );
  AOI2BB2XL U78 ( .B0(addr[5]), .B1(n101), .A0N(n15), .A1N(n112), .Y(n110) );
  OAI211X1 U79 ( .A0(n2), .A1(n147), .B0(n146), .C0(n145), .Y(dout[4]) );
  AOI222XL U80 ( .A0(n144), .A1(n85), .B0(n143), .B1(n142), .C0(n141), .C1(n18), .Y(n145) );
  OA22X1 U81 ( .A0(n81), .A1(n137), .B0(n136), .B1(n18), .Y(n146) );
  NAND3X1 U82 ( .A(n129), .B(n128), .C(n127), .Y(dout[3]) );
  AOI32XL U83 ( .A0(n120), .A1(n85), .A2(addr[1]), .B0(n119), .B1(n118), .Y(
        n128) );
  AOI222XL U84 ( .A0(n144), .A1(n83), .B0(n126), .B1(n16), .C0(n125), .C1(n124), .Y(n127) );
  NAND3BX1 U85 ( .AN(n95), .B(n94), .C(n93), .Y(dout[1]) );
  OAI222X1 U86 ( .A0(n140), .A1(n4), .B0(n112), .B1(n15), .C0(n8), .C1(n91), 
        .Y(n95) );
  AOI32XL U87 ( .A0(addr[1]), .A1(n18), .A2(n125), .B0(n130), .B1(n92), .Y(n93) );
  CLKINVX3 U88 ( .A(n5), .Y(n15) );
  CLKINVX3 U89 ( .A(addr[6]), .Y(n17) );
endmodule


module sbox7_9 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148;

  OAI222X4 U19 ( .A0(n86), .A1(n129), .B0(n4), .B1(n18), .C0(addr[1]), .C1(n8), 
        .Y(n122) );
  OAI33X4 U33 ( .A0(addr[1]), .A1(n4), .A2(n5), .B0(n84), .B1(n6), .B2(n14), 
        .Y(n97) );
  NOR2X2 U44 ( .A(n17), .B(n4), .Y(n116) );
  NOR2X2 U48 ( .A(addr[1]), .B(addr[6]), .Y(n136) );
  NOR2X2 U51 ( .A(n20), .B(n17), .Y(n125) );
  NOR2X2 U52 ( .A(n84), .B(addr[3]), .Y(n131) );
  NOR2X2 U58 ( .A(n93), .B(n124), .Y(n142) );
  NOR2X2 U60 ( .A(n85), .B(addr[1]), .Y(n93) );
  NOR2X2 U62 ( .A(n12), .B(n3), .Y(n137) );
  NOR2X2 U65 ( .A(n85), .B(n87), .Y(n140) );
  NAND2X1 U1 ( .A(n3), .B(n4), .Y(n119) );
  CLKBUFX3 U2 ( .A(addr[4]), .Y(n4) );
  CLKINVX1 U3 ( .A(n12), .Y(n1) );
  CLKINVX1 U4 ( .A(n6), .Y(n2) );
  CLKBUFX3 U5 ( .A(addr[2]), .Y(n5) );
  OAI31X1 U6 ( .A0(n17), .A1(n12), .A2(n87), .B0(n117), .Y(n121) );
  NOR2X4 U7 ( .A(n87), .B(addr[6]), .Y(n124) );
  OAI22X1 U8 ( .A0(addr[1]), .A1(n8), .B0(n5), .B1(n113), .Y(n100) );
  OAI22X1 U9 ( .A0(n4), .A1(n20), .B0(addr[3]), .B1(n11), .Y(n103) );
  AOI211XL U10 ( .A0(n5), .A1(n83), .B0(n131), .C0(n130), .Y(n132) );
  NOR3XL U11 ( .A(n86), .B(addr[3]), .C(n2), .Y(n130) );
  OAI21XL U12 ( .A0(n3), .A1(n1), .B0(n119), .Y(n89) );
  BUFX4 U13 ( .A(addr[5]), .Y(n3) );
  AOI221XL U14 ( .A0(n140), .A1(n89), .B0(n109), .B1(n83), .C0(n88), .Y(n96)
         );
  CLKINVX1 U15 ( .A(n140), .Y(n84) );
  OAI2BB2XL U16 ( .B0(n142), .B1(n11), .A0N(n141), .A1N(n140), .Y(n143) );
  CLKINVX1 U17 ( .A(n125), .Y(n16) );
  CLKINVX1 U18 ( .A(n142), .Y(n83) );
  NAND2X1 U20 ( .A(n16), .B(n19), .Y(n105) );
  CLKINVX1 U21 ( .A(n123), .Y(n7) );
  CLKINVX1 U22 ( .A(n109), .Y(n10) );
  NAND2X1 U23 ( .A(n124), .B(n17), .Y(n113) );
  CLKINVX1 U24 ( .A(n137), .Y(n11) );
  NOR2X1 U25 ( .A(n11), .B(n17), .Y(n109) );
  CLKINVX1 U26 ( .A(n136), .Y(n86) );
  OAI22XL U27 ( .A0(n137), .A1(n18), .B0(n87), .B1(n10), .Y(n146) );
  OAI21X1 U28 ( .A0(n12), .A1(n16), .B0(n129), .Y(n141) );
  NAND2X1 U29 ( .A(n116), .B(n20), .Y(n129) );
  CLKINVX1 U30 ( .A(n93), .Y(n21) );
  OAI21XL U31 ( .A0(n119), .A1(n21), .B0(n118), .Y(n120) );
  OAI21XL U32 ( .A0(n125), .A1(n137), .B0(n124), .Y(n118) );
  NOR2X1 U34 ( .A(n20), .B(n8), .Y(n123) );
  CLKINVX1 U35 ( .A(n145), .Y(n8) );
  OAI22XL U36 ( .A0(n137), .A1(n113), .B0(n85), .B1(n7), .Y(n88) );
  CLKINVX1 U37 ( .A(n116), .Y(n14) );
  CLKINVX1 U38 ( .A(n131), .Y(n18) );
  CLKINVX1 U39 ( .A(n134), .Y(n19) );
  NOR2XL U40 ( .A(n125), .B(n12), .Y(n110) );
  CLKINVX1 U41 ( .A(n119), .Y(n13) );
  CLKINVX1 U42 ( .A(n103), .Y(n9) );
  OA21XL U43 ( .A0(n15), .A1(n21), .B0(n117), .Y(n102) );
  CLKINVX1 U45 ( .A(n105), .Y(n15) );
  OAI2BB1XL U46 ( .A0N(n103), .A1N(n124), .B0(n102), .Y(n104) );
  OAI22X1 U47 ( .A0(n20), .A1(n14), .B0(n4), .B1(n19), .Y(n112) );
  NOR4X1 U49 ( .A(n4), .B(addr[3]), .C(n87), .D(n6), .Y(n99) );
  XNOR2X1 U50 ( .A(addr[6]), .B(n5), .Y(n101) );
  AOI211X1 U53 ( .A0(n116), .A1(addr[6]), .B0(n115), .C0(n114), .Y(n128) );
  OAI222X1 U54 ( .A0(n111), .A1(n84), .B0(n110), .B1(n21), .C0(n86), .C1(n10), 
        .Y(n115) );
  OAI2BB2XL U55 ( .B0(n13), .B1(n113), .A0N(n87), .A1N(n112), .Y(n114) );
  OA21XL U56 ( .A0(n17), .A1(n3), .B0(n7), .Y(n111) );
  NAND2X1 U57 ( .A(n5), .B(n136), .Y(n133) );
  CLKINVX1 U59 ( .A(addr[6]), .Y(n85) );
  AOI211X1 U61 ( .A0(n131), .A1(n3), .B0(n92), .C0(n91), .Y(n95) );
  OAI221X1 U63 ( .A0(n87), .A1(n8), .B0(n84), .B1(n11), .C0(n102), .Y(n92) );
  OAI31X1 U64 ( .A0(n17), .A1(n12), .A2(n86), .B0(n90), .Y(n91) );
  AO21XL U66 ( .A0(n119), .A1(n129), .B0(addr[6]), .Y(n90) );
  NOR2X1 U67 ( .A(n12), .B(addr[3]), .Y(n145) );
  AOI21XL U68 ( .A0(addr[3]), .A1(n98), .B0(n97), .Y(n108) );
  OAI2BB1XL U69 ( .A0N(n6), .A1N(n124), .B0(n133), .Y(n98) );
  NAND3X1 U70 ( .A(n136), .B(n17), .C(n3), .Y(n117) );
  NOR2X1 U71 ( .A(addr[3]), .B(n3), .Y(n134) );
  OAI21X1 U72 ( .A0(n5), .A1(n142), .B0(n133), .Y(n138) );
  OAI22XL U73 ( .A0(n142), .A1(n14), .B0(n1), .B1(n132), .Y(n135) );
  AO21X1 U74 ( .A0(n139), .A1(n20), .B0(n138), .Y(n144) );
  OAI21XL U75 ( .A0(n2), .A1(n87), .B0(n21), .Y(n139) );
  OAI221X1 U76 ( .A0(n96), .A1(n6), .B0(n5), .B1(n95), .C0(n94), .Y(dout[1])
         );
  AOI2BB2X1 U77 ( .B0(n93), .B1(n112), .A0N(n133), .A1N(n9), .Y(n94) );
  OAI211X1 U78 ( .A0(n128), .A1(n6), .B0(n127), .C0(n126), .Y(dout[3]) );
  AOI32XL U79 ( .A0(n125), .A1(n1), .A2(n124), .B0(n123), .B1(n136), .Y(n126)
         );
  OAI31X1 U80 ( .A0(n122), .A1(n121), .A2(n120), .B0(n6), .Y(n127) );
  OAI221X1 U81 ( .A0(n3), .A1(n108), .B0(n107), .B1(n20), .C0(n106), .Y(
        dout[2]) );
  AOI32XL U82 ( .A0(n105), .A1(n6), .A2(n140), .B0(n2), .B1(n104), .Y(n106) );
  AOI211X1 U83 ( .A0(n101), .A1(n4), .B0(n100), .C0(n99), .Y(n107) );
  NAND2X1 U84 ( .A(n148), .B(n147), .Y(dout[4]) );
  AOI222XL U85 ( .A0(n136), .A1(n141), .B0(n3), .B1(n135), .C0(n134), .C1(n138), .Y(n148) );
  AOI222XL U86 ( .A0(n5), .A1(n146), .B0(n145), .B1(n144), .C0(n143), .C1(n6), 
        .Y(n147) );
  CLKINVX3 U87 ( .A(n5), .Y(n6) );
  CLKINVX3 U88 ( .A(n4), .Y(n12) );
  CLKINVX3 U89 ( .A(addr[3]), .Y(n17) );
  CLKINVX3 U90 ( .A(n3), .Y(n20) );
  CLKINVX3 U91 ( .A(addr[1]), .Y(n87) );
endmodule


module sbox8_9 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132;

  NAND2X2 U41 ( .A(addr[6]), .B(n15), .Y(n131) );
  NAND2X2 U48 ( .A(addr[4]), .B(n11), .Y(n123) );
  NAND2X2 U49 ( .A(n2), .B(n12), .Y(n87) );
  NAND2X2 U50 ( .A(addr[1]), .B(n75), .Y(n124) );
  NAND2X2 U54 ( .A(addr[2]), .B(n9), .Y(n116) );
  NAND2X2 U60 ( .A(addr[6]), .B(addr[1]), .Y(n105) );
  NAND2X2 U61 ( .A(n15), .B(n75), .Y(n108) );
  OAI31X1 U1 ( .A0(n123), .A1(addr[6]), .A2(n116), .B0(n109), .Y(n110) );
  AOI222X1 U2 ( .A0(n88), .A1(addr[2]), .B0(n12), .B1(n4), .C0(n5), .C1(n92), 
        .Y(n114) );
  OAI222X1 U3 ( .A0(addr[2]), .A1(n126), .B0(n11), .B1(n125), .C0(n124), .C1(
        n123), .Y(n127) );
  NAND2X4 U4 ( .A(addr[4]), .B(n2), .Y(n115) );
  OAI32X1 U5 ( .A0(n75), .A1(addr[4]), .A2(n92), .B0(n115), .B1(n108), .Y(n96)
         );
  OAI221X1 U6 ( .A0(n105), .A1(n87), .B0(addr[4]), .B1(n108), .C0(n86), .Y(n90) );
  AOI32XL U7 ( .A0(n74), .A1(n7), .A2(n2), .B0(n14), .B1(n117), .Y(n130) );
  OA21XL U8 ( .A0(n5), .A1(n9), .B0(n121), .Y(n78) );
  INVXL U9 ( .A(n119), .Y(n3) );
  INVX3 U10 ( .A(n2), .Y(n11) );
  BUFX4 U11 ( .A(addr[3]), .Y(n2) );
  CLKBUFX3 U12 ( .A(addr[5]), .Y(n1) );
  CLKINVX1 U13 ( .A(n108), .Y(n14) );
  CLKINVX1 U14 ( .A(n107), .Y(n6) );
  CLKINVX1 U15 ( .A(n93), .Y(n10) );
  NAND2X1 U16 ( .A(n11), .B(n12), .Y(n93) );
  NAND2X1 U17 ( .A(n5), .B(n9), .Y(n121) );
  OAI21XL U18 ( .A0(n115), .A1(n9), .B0(n107), .Y(n77) );
  OAI21X1 U19 ( .A0(n12), .A1(n9), .B0(n123), .Y(n88) );
  OAI31XL U20 ( .A0(n115), .A1(n15), .A2(n116), .B0(n118), .Y(n94) );
  CLKINVX1 U21 ( .A(n131), .Y(n13) );
  NAND2X1 U22 ( .A(n7), .B(n11), .Y(n107) );
  OAI22XL U23 ( .A0(n116), .A1(n123), .B0(n7), .B1(n115), .Y(n117) );
  OAI22XL U24 ( .A0(n123), .A1(n108), .B0(n131), .B1(n93), .Y(n95) );
  OAI2BB2XL U25 ( .B0(n115), .B1(n131), .A0N(n88), .A1N(n16), .Y(n89) );
  AOI211XL U26 ( .A0(n108), .A1(n105), .B0(n12), .C0(n121), .Y(n85) );
  CLKINVX1 U27 ( .A(n124), .Y(n74) );
  OAI22XL U28 ( .A0(n7), .A1(n123), .B0(n78), .B1(n87), .Y(n81) );
  NAND2BX2 U29 ( .AN(n78), .B(n11), .Y(n120) );
  NAND2XL U30 ( .A(n115), .B(n93), .Y(n104) );
  OAI2BB2XL U31 ( .B0(n106), .B1(n105), .A0N(n104), .A1N(n74), .Y(n111) );
  NOR2BXL U32 ( .AN(n123), .B(n103), .Y(n106) );
  NAND3X1 U33 ( .A(n104), .B(n15), .C(n7), .Y(n84) );
  AO21X1 U34 ( .A0(n7), .A1(n16), .B0(n101), .Y(n102) );
  OAI33X1 U35 ( .A0(n75), .A1(n11), .A2(n100), .B0(n5), .B1(n103), .B2(n124), 
        .Y(n101) );
  OA22XL U36 ( .A0(n107), .A1(n131), .B0(n120), .B1(n124), .Y(n98) );
  CLKINVX1 U37 ( .A(n125), .Y(n8) );
  OAI21XL U38 ( .A0(n74), .A1(n13), .B0(addr[4]), .Y(n86) );
  NAND2X1 U39 ( .A(n1), .B(n5), .Y(n100) );
  OAI221X1 U40 ( .A0(n124), .A1(n121), .B0(addr[1]), .B1(n120), .C0(n3), .Y(
        n128) );
  OAI31XL U42 ( .A0(n5), .A1(n15), .A2(n11), .B0(n118), .Y(n119) );
  NAND2X1 U43 ( .A(n16), .B(addr[2]), .Y(n125) );
  NAND4XL U44 ( .A(n13), .B(n1), .C(n2), .D(addr[2]), .Y(n109) );
  NAND3X1 U45 ( .A(n7), .B(n75), .C(n2), .Y(n118) );
  OAI21XL U46 ( .A0(n1), .A1(n87), .B0(n114), .Y(n76) );
  OAI22XL U47 ( .A0(n108), .A1(n120), .B0(n79), .B1(n100), .Y(n80) );
  AOI221XL U51 ( .A0(n13), .A1(n11), .B0(n16), .B1(n2), .C0(n91), .Y(n79) );
  NOR2X1 U52 ( .A(n1), .B(n2), .Y(n103) );
  NOR2X1 U53 ( .A(n87), .B(addr[6]), .Y(n91) );
  NOR2X1 U55 ( .A(n11), .B(n1), .Y(n92) );
  CLKINVX1 U56 ( .A(n100), .Y(n4) );
  OA21XL U57 ( .A0(n1), .A1(n115), .B0(n120), .Y(n132) );
  AOI221XL U58 ( .A0(n14), .A1(n2), .B0(n16), .B1(addr[4]), .C0(n122), .Y(n126) );
  OAI22XL U59 ( .A0(n2), .A1(n15), .B0(addr[4]), .B1(n131), .Y(n122) );
  OAI211X1 U62 ( .A0(addr[2]), .A1(n99), .B0(n98), .C0(n97), .Y(dout[2]) );
  AOI221XL U63 ( .A0(addr[2]), .A1(n96), .B0(n1), .B1(n95), .C0(n94), .Y(n97)
         );
  AOI221XL U64 ( .A0(n91), .A1(n1), .B0(n90), .B1(n9), .C0(n89), .Y(n99) );
  OAI211X1 U65 ( .A0(n132), .A1(n131), .B0(n130), .C0(n129), .Y(dout[4]) );
  AOI222XL U66 ( .A0(n128), .A1(n12), .B0(n1), .B1(n127), .C0(n6), .C1(n16), 
        .Y(n129) );
  OAI211X1 U67 ( .A0(addr[1]), .A1(n114), .B0(n113), .C0(n112), .Y(dout[3]) );
  AOI221XL U68 ( .A0(n111), .A1(n5), .B0(n6), .B1(n14), .C0(n110), .Y(n112) );
  AOI2BB2XL U69 ( .B0(n102), .B1(n12), .A0N(n115), .A1N(n125), .Y(n113) );
  NAND4BX1 U70 ( .AN(n85), .B(n84), .C(n83), .D(n82), .Y(dout[1]) );
  AOI221XL U71 ( .A0(n13), .A1(n81), .B0(n10), .B1(n8), .C0(n80), .Y(n82) );
  AOI22X1 U72 ( .A0(n16), .A1(n77), .B0(n74), .B1(n76), .Y(n83) );
  CLKINVX3 U73 ( .A(addr[2]), .Y(n5) );
  CLKINVX3 U74 ( .A(n116), .Y(n7) );
  CLKINVX3 U75 ( .A(n1), .Y(n9) );
  CLKINVX3 U76 ( .A(addr[4]), .Y(n12) );
  CLKINVX3 U77 ( .A(addr[1]), .Y(n15) );
  CLKINVX3 U78 ( .A(n105), .Y(n16) );
  CLKINVX3 U79 ( .A(addr[6]), .Y(n75) );
endmodule


module crp_9 ( P, R, K_sub );
  output [1:32] P;
  input [1:32] R;
  input [1:48] K_sub;
  wire   n1;
  wire   [1:48] X;

  sbox1_9 u0 ( .addr(X[1:6]), .dout({P[9], P[17], P[23], P[31]}) );
  sbox2_9 u1 ( .addr({X[7], n1, X[9:12]}), .dout({P[13], P[28], P[2], P[18]})
         );
  sbox3_9 u2 ( .addr(X[13:18]), .dout({P[24], P[16], P[30], P[6]}) );
  sbox4_9 u3 ( .addr(X[19:24]), .dout({P[26], P[20], P[10], P[1]}) );
  sbox5_9 u4 ( .addr(X[25:30]), .dout({P[8], P[14], P[25], P[3]}) );
  sbox6_9 u5 ( .addr(X[31:36]), .dout({P[4], P[29], P[11], P[19]}) );
  sbox7_9 u6 ( .addr(X[37:42]), .dout({P[32], P[12], P[22], P[7]}) );
  sbox8_9 u7 ( .addr(X[43:48]), .dout({P[5], P[27], P[15], P[21]}) );
  XOR2X1 U1 ( .A(R[1]), .B(K_sub[2]), .Y(X[2]) );
  CLKXOR2X4 U2 ( .A(R[29]), .B(K_sub[42]), .Y(X[42]) );
  CLKXOR2X4 U3 ( .A(R[5]), .B(K_sub[6]), .Y(X[6]) );
  CLKXOR2X4 U4 ( .A(R[16]), .B(K_sub[25]), .Y(X[25]) );
  CLKXOR2X4 U5 ( .A(R[22]), .B(K_sub[33]), .Y(X[33]) );
  CLKXOR2X4 U6 ( .A(R[8]), .B(K_sub[11]), .Y(X[11]) );
  CLKXOR2X4 U7 ( .A(R[29]), .B(K_sub[44]), .Y(X[44]) );
  CLKXOR2X4 U8 ( .A(R[12]), .B(K_sub[19]), .Y(X[19]) );
  CLKXOR2X4 U9 ( .A(R[10]), .B(K_sub[15]), .Y(X[15]) );
  XNOR2X1 U10 ( .A(R[5]), .B(K_sub[8]), .Y(X[8]) );
  INVX3 U11 ( .A(X[8]), .Y(n1) );
  CLKXOR2X4 U12 ( .A(R[20]), .B(K_sub[31]), .Y(X[31]) );
  CLKXOR2X4 U13 ( .A(R[16]), .B(K_sub[23]), .Y(X[23]) );
  CLKXOR2X4 U14 ( .A(R[31]), .B(K_sub[46]), .Y(X[46]) );
  CLKXOR2X4 U15 ( .A(R[26]), .B(K_sub[39]), .Y(X[39]) );
  CLKXOR2X4 U16 ( .A(R[20]), .B(K_sub[29]), .Y(X[29]) );
  CLKXOR2X2 U17 ( .A(R[4]), .B(K_sub[5]), .Y(X[5]) );
  CLKXOR2X2 U18 ( .A(R[15]), .B(K_sub[22]), .Y(X[22]) );
  CLKXOR2X2 U19 ( .A(R[24]), .B(K_sub[35]), .Y(X[35]) );
  CLKXOR2X2 U20 ( .A(R[21]), .B(K_sub[30]), .Y(X[30]) );
  CLKXOR2X2 U21 ( .A(R[12]), .B(K_sub[17]), .Y(X[17]) );
  CLKXOR2X2 U22 ( .A(R[32]), .B(K_sub[1]), .Y(X[1]) );
  CLKXOR2X2 U23 ( .A(R[13]), .B(K_sub[20]), .Y(X[20]) );
  CLKXOR2X2 U24 ( .A(R[18]), .B(K_sub[27]), .Y(X[27]) );
  CLKXOR2X2 U25 ( .A(R[8]), .B(K_sub[13]), .Y(X[13]) );
  CLKXOR2X2 U26 ( .A(R[4]), .B(K_sub[7]), .Y(X[7]) );
  CLKXOR2X2 U27 ( .A(R[24]), .B(K_sub[37]), .Y(X[37]) );
  CLKXOR2X2 U28 ( .A(R[28]), .B(K_sub[43]), .Y(X[43]) );
  CLKXOR2X2 U29 ( .A(R[1]), .B(K_sub[48]), .Y(X[48]) );
  CLKXOR2X2 U30 ( .A(R[17]), .B(K_sub[24]), .Y(X[24]) );
  CLKXOR2X2 U31 ( .A(R[9]), .B(K_sub[12]), .Y(X[12]) );
  CLKXOR2X2 U32 ( .A(R[13]), .B(K_sub[18]), .Y(X[18]) );
  CLKXOR2X2 U33 ( .A(R[25]), .B(K_sub[36]), .Y(X[36]) );
  XOR2X1 U34 ( .A(R[23]), .B(K_sub[34]), .Y(X[34]) );
  XOR2X1 U35 ( .A(R[9]), .B(K_sub[14]), .Y(X[14]) );
  XOR2X1 U36 ( .A(R[30]), .B(K_sub[45]), .Y(X[45]) );
  XOR2X1 U37 ( .A(R[21]), .B(K_sub[32]), .Y(X[32]) );
  XOR2X1 U38 ( .A(R[25]), .B(K_sub[38]), .Y(X[38]) );
  XOR2X1 U39 ( .A(R[27]), .B(K_sub[40]), .Y(X[40]) );
  XOR2X1 U40 ( .A(R[3]), .B(K_sub[4]), .Y(X[4]) );
  XOR2X1 U41 ( .A(R[11]), .B(K_sub[16]), .Y(X[16]) );
  XOR2X1 U42 ( .A(R[7]), .B(K_sub[10]), .Y(X[10]) );
  XOR2X1 U43 ( .A(R[14]), .B(K_sub[21]), .Y(X[21]) );
  XOR2X1 U44 ( .A(R[6]), .B(K_sub[9]), .Y(X[9]) );
  XOR2X1 U45 ( .A(R[2]), .B(K_sub[3]), .Y(X[3]) );
  XOR2X1 U46 ( .A(R[28]), .B(K_sub[41]), .Y(X[41]) );
  XOR2X1 U47 ( .A(R[17]), .B(K_sub[26]), .Y(X[26]) );
  XOR2X1 U48 ( .A(R[32]), .B(K_sub[47]), .Y(X[47]) );
  XOR2X1 U49 ( .A(R[19]), .B(K_sub[28]), .Y(X[28]) );
endmodule


module sbox1_8 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127;

  OAI222X4 U13 ( .A0(addr[5]), .A1(n101), .B0(n1), .B1(n100), .C0(n99), .C1(n8), .Y(dout[3]) );
  OAI21X2 U42 ( .A0(n4), .A1(n112), .B0(n106), .Y(n123) );
  NAND2X2 U44 ( .A(addr[6]), .B(n70), .Y(n115) );
  NAND2X2 U48 ( .A(addr[1]), .B(n11), .Y(n114) );
  OAI22X2 U49 ( .A0(n71), .A1(n6), .B0(addr[5]), .B1(n120), .Y(n85) );
  NAND2X2 U50 ( .A(n3), .B(n71), .Y(n120) );
  NOR2X2 U51 ( .A(n71), .B(n3), .Y(n124) );
  NOR3X2 U55 ( .A(n2), .B(addr[6]), .C(n8), .Y(n102) );
  NOR2X2 U56 ( .A(n109), .B(n3), .Y(n93) );
  NAND2X2 U57 ( .A(addr[1]), .B(addr[6]), .Y(n109) );
  NAND2X2 U59 ( .A(n70), .B(n11), .Y(n112) );
  NOR2X1 U1 ( .A(n114), .B(n120), .Y(n104) );
  BUFX4 U2 ( .A(addr[4]), .Y(n2) );
  CLKBUFX3 U3 ( .A(addr[2]), .Y(n1) );
  OAI32X1 U4 ( .A0(n112), .A1(n2), .A2(n4), .B0(n115), .B1(n113), .Y(n80) );
  NOR2BXL U5 ( .AN(n118), .B(n1), .Y(n122) );
  CLKBUFX3 U6 ( .A(addr[2]), .Y(n4) );
  INVX3 U7 ( .A(addr[6]), .Y(n11) );
  OAI221X4 U8 ( .A0(n88), .A1(n6), .B0(addr[5]), .B1(n87), .C0(n86), .Y(
        dout[2]) );
  OAI221X4 U9 ( .A0(addr[5]), .A1(n127), .B0(n126), .B1(n6), .C0(n125), .Y(
        dout[4]) );
  OA21XL U10 ( .A0(n95), .A1(n115), .B0(n107), .Y(n119) );
  AOI222XL U11 ( .A0(n10), .A1(n1), .B0(n2), .B1(n110), .C0(n12), .C1(n8), .Y(
        n111) );
  AOI2BB2X1 U12 ( .B0(n2), .B1(n12), .A0N(addr[4]), .A1N(n115), .Y(n91) );
  BUFX4 U14 ( .A(addr[3]), .Y(n3) );
  CLKINVX1 U15 ( .A(n112), .Y(n10) );
  CLKINVX1 U16 ( .A(n113), .Y(n7) );
  NAND2BX1 U17 ( .AN(n104), .B(n119), .Y(n84) );
  CLKXOR2X2 U18 ( .A(n72), .B(n8), .Y(n90) );
  NOR2X1 U19 ( .A(n71), .B(n72), .Y(n118) );
  OAI21XL U20 ( .A0(n72), .A1(n114), .B0(n91), .Y(n92) );
  NAND2X1 U21 ( .A(n93), .B(n71), .Y(n107) );
  NAND2X1 U22 ( .A(n8), .B(n72), .Y(n113) );
  OAI211X1 U23 ( .A0(n71), .A1(n114), .B0(n108), .C0(n107), .Y(n89) );
  CLKINVX1 U24 ( .A(n109), .Y(n12) );
  NAND2X1 U25 ( .A(n124), .B(n69), .Y(n108) );
  CLKINVX1 U26 ( .A(n114), .Y(n9) );
  CLKINVX1 U27 ( .A(n115), .Y(n69) );
  CLKINVX1 U28 ( .A(n95), .Y(n5) );
  AO22X1 U29 ( .A0(n90), .A1(n69), .B0(n72), .B1(n123), .Y(n76) );
  OAI31X1 U30 ( .A0(n8), .A1(n3), .A2(n70), .B0(n103), .Y(n105) );
  AOI31XL U31 ( .A0(n70), .A1(n8), .A2(n2), .B0(n102), .Y(n103) );
  AOI211X1 U32 ( .A0(n13), .A1(n4), .B0(n117), .C0(n116), .Y(n126) );
  CLKINVX1 U33 ( .A(n108), .Y(n13) );
  AOI211X1 U34 ( .A0(n115), .A1(n114), .B0(n113), .C0(n2), .Y(n116) );
  OAI22X1 U35 ( .A0(n120), .A1(n112), .B0(n111), .B1(n72), .Y(n117) );
  AOI211X1 U36 ( .A0(n12), .A1(n118), .B0(n81), .C0(n80), .Y(n88) );
  OAI22X1 U37 ( .A0(n91), .A1(n8), .B0(n3), .B1(n106), .Y(n81) );
  CLKINVX3 U38 ( .A(addr[5]), .Y(n6) );
  NAND2X1 U39 ( .A(n3), .B(n6), .Y(n95) );
  NAND2X1 U40 ( .A(n9), .B(n1), .Y(n106) );
  XOR2X1 U41 ( .A(n82), .B(n2), .Y(n83) );
  NAND2X1 U43 ( .A(n1), .B(n3), .Y(n82) );
  OAI22XL U45 ( .A0(n3), .A1(n70), .B0(n72), .B1(n112), .Y(n94) );
  AOI211XL U46 ( .A0(n98), .A1(n72), .B0(n97), .C0(n104), .Y(n99) );
  OAI22XL U47 ( .A0(n96), .A1(n71), .B0(n95), .B1(n109), .Y(n97) );
  OAI22XL U52 ( .A0(n11), .A1(n6), .B0(n2), .B1(addr[1]), .Y(n98) );
  AOI221XL U53 ( .A0(n5), .A1(addr[6]), .B0(addr[5]), .B1(n94), .C0(n93), .Y(
        n96) );
  OAI21XL U54 ( .A0(addr[1]), .A1(n120), .B0(n119), .Y(n121) );
  AOI221XL U58 ( .A0(n10), .A1(n118), .B0(n93), .B1(n6), .C0(n75), .Y(n78) );
  OAI31X1 U60 ( .A0(n6), .A1(n2), .A2(n74), .B0(n73), .Y(n75) );
  OA21XL U61 ( .A0(n3), .A1(n11), .B0(n109), .Y(n74) );
  OAI21XL U62 ( .A0(n124), .A1(n85), .B0(n9), .Y(n73) );
  OAI21XL U63 ( .A0(n1), .A1(n70), .B0(n109), .Y(n110) );
  INVX4 U64 ( .A(n4), .Y(n8) );
  AOI222XL U65 ( .A0(n124), .A1(n123), .B0(n122), .B1(addr[6]), .C0(n1), .C1(
        n121), .Y(n125) );
  NOR4BBX1 U66 ( .AN(n107), .BN(n106), .C(n105), .D(n104), .Y(n127) );
  AOI222XL U67 ( .A0(n10), .A1(n90), .B0(n89), .B1(n8), .C0(n123), .C1(n71), 
        .Y(n101) );
  AOI2BB2XL U68 ( .B0(addr[5]), .B1(n92), .A0N(n120), .A1N(addr[1]), .Y(n100)
         );
  AOI32X1 U69 ( .A0(n4), .A1(n85), .A2(n10), .B0(n84), .B1(n8), .Y(n86) );
  AOI222XL U70 ( .A0(n124), .A1(n70), .B0(n83), .B1(addr[1]), .C0(n7), .C1(n11), .Y(n87) );
  OAI221X1 U71 ( .A0(n79), .A1(n6), .B0(n4), .B1(n78), .C0(n77), .Y(dout[1])
         );
  AOI32XL U72 ( .A0(addr[6]), .A1(n85), .A2(n1), .B0(n76), .B1(n6), .Y(n77) );
  AOI221X1 U73 ( .A0(n10), .A1(n90), .B0(n4), .B1(n93), .C0(n102), .Y(n79) );
  CLKINVX3 U74 ( .A(addr[1]), .Y(n70) );
  CLKINVX3 U75 ( .A(n2), .Y(n71) );
  CLKINVX3 U76 ( .A(n3), .Y(n72) );
endmodule


module sbox2_8 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147;

  NAND2X2 U55 ( .A(n2), .B(n82), .Y(n136) );
  NAND2X2 U57 ( .A(addr[2]), .B(n5), .Y(n104) );
  NAND2X2 U60 ( .A(addr[5]), .B(addr[2]), .Y(n132) );
  NOR2X2 U61 ( .A(n10), .B(n8), .Y(n101) );
  NAND2X2 U62 ( .A(n83), .B(n9), .Y(n146) );
  NAND2X2 U63 ( .A(n3), .B(n13), .Y(n124) );
  NAND2X2 U64 ( .A(addr[6]), .B(n83), .Y(n122) );
  NAND2X2 U67 ( .A(n3), .B(n2), .Y(n133) );
  AOI222XL U1 ( .A0(n14), .A1(n7), .B0(n88), .B1(n13), .C0(n140), .C1(n8), .Y(
        n89) );
  CLKINVX1 U2 ( .A(n121), .Y(n10) );
  AOI211X1 U3 ( .A0(n6), .A1(n95), .B0(n94), .C0(n93), .Y(n96) );
  NOR2X1 U4 ( .A(n104), .B(n2), .Y(n141) );
  NOR2X1 U5 ( .A(n124), .B(n2), .Y(n140) );
  CLKBUFX4 U6 ( .A(addr[4]), .Y(n2) );
  CLKINVX1 U7 ( .A(addr[5]), .Y(n1) );
  OAI22X1 U8 ( .A0(n117), .A1(n114), .B0(n89), .B1(n5), .Y(n94) );
  INVX3 U9 ( .A(addr[5]), .Y(n5) );
  OAI211X4 U10 ( .A0(n147), .A1(n146), .B0(n145), .C0(n144), .Y(dout[4]) );
  NAND2X1 U11 ( .A(addr[1]), .B(addr[6]), .Y(n121) );
  CLKINVX2 U12 ( .A(addr[1]), .Y(n83) );
  OAI221X1 U13 ( .A0(addr[1]), .A1(n136), .B0(n133), .B1(n83), .C0(n87), .Y(
        n95) );
  NAND2X4 U14 ( .A(addr[1]), .B(n9), .Y(n114) );
  INVX3 U15 ( .A(addr[6]), .Y(n9) );
  NAND2XL U16 ( .A(n102), .B(n82), .Y(n109) );
  AOI2BB2X1 U17 ( .B0(n5), .B1(n12), .A0N(n104), .A1N(n136), .Y(n117) );
  NOR3BXL U18 ( .AN(n135), .B(n134), .C(n14), .Y(n147) );
  BUFX4 U19 ( .A(addr[3]), .Y(n3) );
  NAND2X1 U20 ( .A(n14), .B(n10), .Y(n113) );
  CLKINVX1 U21 ( .A(n146), .Y(n8) );
  CLKINVX1 U22 ( .A(n115), .Y(n14) );
  CLKINVX1 U23 ( .A(n122), .Y(n11) );
  OAI31X1 U24 ( .A0(n124), .A1(n9), .A2(n5), .B0(n123), .Y(n128) );
  OAI21XL U25 ( .A0(n1), .A1(n83), .B0(n140), .Y(n123) );
  OAI22X1 U26 ( .A0(n122), .A1(n124), .B0(n101), .B1(n132), .Y(n84) );
  INVX1 U27 ( .A(n114), .Y(n7) );
  OAI22X1 U28 ( .A0(n122), .A1(n82), .B0(n15), .B1(n121), .Y(n129) );
  NAND3X1 U29 ( .A(n15), .B(n5), .C(n83), .Y(n111) );
  NAND2X1 U30 ( .A(n82), .B(n15), .Y(n115) );
  OAI21XL U31 ( .A0(n13), .A1(n133), .B0(n135), .Y(n85) );
  OAI22XL U32 ( .A0(n117), .A1(n146), .B0(n116), .B1(n132), .Y(n118) );
  AOI222XL U33 ( .A0(n7), .A1(n115), .B0(n16), .B1(n9), .C0(n14), .C1(n8), .Y(
        n116) );
  CLKINVX1 U34 ( .A(n104), .Y(n4) );
  OAI2BB2XL U35 ( .B0(n114), .B1(n135), .A0N(n126), .A1N(n16), .Y(n106) );
  OAI21XL U36 ( .A0(n112), .A1(n114), .B0(n111), .Y(n120) );
  OAI21XL U37 ( .A0(n133), .A1(n114), .B0(n113), .Y(n119) );
  CLKINVX1 U38 ( .A(n124), .Y(n12) );
  CLKINVX1 U39 ( .A(n136), .Y(n81) );
  CLKINVX1 U40 ( .A(n133), .Y(n16) );
  CLKINVX1 U41 ( .A(n132), .Y(n6) );
  AOI2BB1X1 U42 ( .A0N(n126), .A1N(n125), .B0(n136), .Y(n127) );
  OAI22XL U43 ( .A0(n104), .A1(n114), .B0(n101), .B1(n132), .Y(n102) );
  AO21XL U44 ( .A0(n13), .A1(n81), .B0(n141), .Y(n86) );
  AO21X1 U45 ( .A0(n82), .A1(n4), .B0(n140), .Y(n142) );
  NAND3X1 U46 ( .A(n13), .B(n15), .C(addr[5]), .Y(n135) );
  OAI22X1 U47 ( .A0(addr[5]), .A1(n121), .B0(n122), .B1(n5), .Y(n126) );
  AOI2BB1X1 U48 ( .A0N(n3), .A1N(n1), .B0(n81), .Y(n112) );
  NOR3X1 U49 ( .A(addr[1]), .B(addr[2]), .C(n5), .Y(n125) );
  AOI2BB1XL U50 ( .A0N(n92), .A1N(n91), .B0(addr[5]), .Y(n93) );
  OAI31XL U51 ( .A0(n114), .A1(n2), .A2(n82), .B0(n90), .Y(n91) );
  OAI21XL U52 ( .A0(n16), .A1(n12), .B0(n11), .Y(n90) );
  NAND2X1 U53 ( .A(n7), .B(n2), .Y(n137) );
  OAI31XL U54 ( .A0(n101), .A1(n3), .A2(addr[2]), .B0(n113), .Y(n92) );
  OAI211X1 U56 ( .A0(n139), .A1(n5), .B0(n138), .C0(n137), .Y(n143) );
  NAND3X1 U58 ( .A(n15), .B(n5), .C(addr[6]), .Y(n138) );
  AOI2BB2X1 U59 ( .B0(n11), .B1(n82), .A0N(n83), .A1N(n136), .Y(n139) );
  OAI22XL U65 ( .A0(addr[5]), .A1(n133), .B0(n3), .B1(n132), .Y(n134) );
  OAI2BB2XL U66 ( .B0(n112), .B1(n122), .A0N(n1), .A1N(n99), .Y(n100) );
  OAI211X1 U68 ( .A0(n146), .A1(n2), .B0(n137), .C0(n113), .Y(n99) );
  NAND3X1 U69 ( .A(n11), .B(n15), .C(n3), .Y(n87) );
  AOI2BB2XL U70 ( .B0(n3), .B1(n105), .A0N(n137), .A1N(n132), .Y(n108) );
  OAI211XL U71 ( .A0(n104), .A1(n146), .B0(n103), .C0(n111), .Y(n105) );
  NAND3XL U72 ( .A(addr[5]), .B(n15), .C(n10), .Y(n103) );
  OAI22XL U73 ( .A0(n3), .A1(n114), .B0(n9), .B1(n115), .Y(n88) );
  NAND4X1 U74 ( .A(n110), .B(n109), .C(n108), .D(n107), .Y(dout[2]) );
  AOI32XL U75 ( .A0(addr[1]), .A1(addr[2]), .A2(n81), .B0(n100), .B1(n13), .Y(
        n110) );
  AOI221XL U76 ( .A0(n125), .A1(addr[4]), .B0(n141), .B1(n11), .C0(n106), .Y(
        n107) );
  AOI33XL U77 ( .A0(n11), .A1(n4), .A2(n2), .B0(n6), .B1(n146), .B2(n3), .Y(
        n145) );
  AOI222XL U78 ( .A0(n143), .A1(n13), .B0(n10), .B1(n142), .C0(n7), .C1(n141), 
        .Y(n144) );
  NAND3X1 U79 ( .A(n98), .B(n97), .C(n96), .Y(dout[1]) );
  AOI32XL U80 ( .A0(n4), .A1(n83), .A2(n14), .B0(n8), .B1(n86), .Y(n97) );
  AOI22X1 U81 ( .A0(n10), .A1(n85), .B0(n2), .B1(n84), .Y(n98) );
  NAND2X1 U82 ( .A(n131), .B(n130), .Y(dout[3]) );
  AOI221XL U83 ( .A0(n120), .A1(n13), .B0(addr[2]), .B1(n119), .C0(n118), .Y(
        n131) );
  AOI211X1 U84 ( .A0(n4), .A1(n129), .B0(n128), .C0(n127), .Y(n130) );
  CLKINVX3 U85 ( .A(addr[2]), .Y(n13) );
  CLKINVX3 U86 ( .A(n2), .Y(n15) );
  CLKINVX3 U87 ( .A(n3), .Y(n82) );
endmodule


module sbox3_8 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134;

  NOR2X2 U35 ( .A(n76), .B(addr[3]), .Y(n109) );
  NOR2X2 U50 ( .A(addr[1]), .B(addr[6]), .Y(n108) );
  NOR2X2 U52 ( .A(n78), .B(n3), .Y(n88) );
  NOR2X2 U56 ( .A(n78), .B(n16), .Y(n95) );
  NOR2X1 U1 ( .A(n76), .B(n78), .Y(n107) );
  OAI221X1 U2 ( .A0(n125), .A1(n76), .B0(n4), .B1(addr[1]), .C0(n14), .Y(n105)
         );
  BUFX4 U3 ( .A(addr[4]), .Y(n3) );
  INVXL U4 ( .A(n2), .Y(n1) );
  NOR2X1 U5 ( .A(n10), .B(n4), .Y(n92) );
  NOR2X1 U6 ( .A(n77), .B(n4), .Y(n122) );
  NOR2X1 U7 ( .A(n14), .B(n4), .Y(n96) );
  NOR2X1 U8 ( .A(n4), .B(n3), .Y(n111) );
  CLKBUFX3 U9 ( .A(addr[2]), .Y(n4) );
  INVX1 U10 ( .A(addr[2]), .Y(n2) );
  OAI33X1 U11 ( .A0(n77), .A1(n126), .A2(n16), .B0(n76), .B1(n95), .B2(n120), 
        .Y(n80) );
  INVX3 U12 ( .A(n4), .Y(n16) );
  OAI221X1 U13 ( .A0(addr[5]), .A1(n91), .B0(n90), .B1(n19), .C0(n89), .Y(
        dout[1]) );
  NOR2X4 U14 ( .A(n11), .B(n79), .Y(n125) );
  NOR2X4 U15 ( .A(addr[3]), .B(n3), .Y(n131) );
  NOR2X4 U16 ( .A(n79), .B(addr[6]), .Y(n126) );
  INVX3 U17 ( .A(addr[1]), .Y(n79) );
  NAND2XL U18 ( .A(n95), .B(n125), .Y(n133) );
  OAI211XL U19 ( .A0(n3), .A1(n9), .B0(n129), .C0(n128), .Y(n130) );
  NAND4XL U20 ( .A(n115), .B(n114), .C(n113), .D(n112), .Y(n116) );
  CLKINVX1 U21 ( .A(n133), .Y(n7) );
  INVX1 U22 ( .A(n125), .Y(n5) );
  CLKINVX1 U23 ( .A(n107), .Y(n20) );
  NAND2X1 U24 ( .A(n10), .B(n12), .Y(n123) );
  CLKINVX1 U25 ( .A(n87), .Y(n12) );
  CLKINVX1 U26 ( .A(n121), .Y(n15) );
  CLKINVX1 U27 ( .A(n120), .Y(n6) );
  CLKINVX1 U28 ( .A(n115), .Y(n8) );
  CLKINVX1 U29 ( .A(n108), .Y(n14) );
  NOR2X1 U30 ( .A(n10), .B(n16), .Y(n104) );
  NOR2X1 U31 ( .A(n5), .B(n16), .Y(n110) );
  INVX1 U32 ( .A(n126), .Y(n13) );
  AOI21X1 U33 ( .A0(n78), .A1(n16), .B0(n95), .Y(n121) );
  OAI21XL U34 ( .A0(n111), .A1(n131), .B0(n125), .Y(n83) );
  CLKINVX1 U36 ( .A(n82), .Y(n10) );
  NOR2X1 U37 ( .A(n13), .B(n76), .Y(n87) );
  NOR2X1 U38 ( .A(n125), .B(n108), .Y(n120) );
  OAI21XL U39 ( .A0(n110), .A1(n92), .B0(n131), .Y(n101) );
  NAND2X1 U40 ( .A(n104), .B(n88), .Y(n115) );
  CLKINVX1 U41 ( .A(n88), .Y(n77) );
  CLKINVX1 U42 ( .A(n92), .Y(n9) );
  CLKINVX1 U43 ( .A(n111), .Y(n17) );
  CLKINVX1 U44 ( .A(n122), .Y(n18) );
  OR2X1 U45 ( .A(n104), .B(n96), .Y(n127) );
  OAI221X1 U46 ( .A0(n13), .A1(n17), .B0(n16), .B1(n12), .C0(n94), .Y(n99) );
  AOI221XL U47 ( .A0(n96), .A1(n3), .B0(n93), .B1(n76), .C0(n7), .Y(n94) );
  OAI21XL U48 ( .A0(n16), .A1(n14), .B0(n9), .Y(n93) );
  XNOR2X1 U49 ( .A(addr[5]), .B(addr[3]), .Y(n103) );
  CLKINVX1 U51 ( .A(addr[5]), .Y(n19) );
  OAI221X1 U53 ( .A0(n14), .A1(n17), .B0(n5), .B1(n77), .C0(n106), .Y(n117) );
  AOI221XL U54 ( .A0(addr[3]), .A1(n105), .B0(n104), .B1(n131), .C0(n7), .Y(
        n106) );
  CLKINVX1 U55 ( .A(addr[6]), .Y(n11) );
  NAND3X1 U57 ( .A(n4), .B(n79), .C(n109), .Y(n114) );
  NOR2X1 U58 ( .A(n11), .B(addr[1]), .Y(n82) );
  AOI32XL U59 ( .A0(n16), .A1(n78), .A2(n125), .B0(n124), .B1(n11), .Y(n129)
         );
  AOI22XL U60 ( .A0(n3), .A1(n127), .B0(n126), .B1(n131), .Y(n128) );
  OAI22XL U61 ( .A0(n3), .A1(n2), .B0(n4), .B1(n20), .Y(n124) );
  AOI222XL U62 ( .A0(n111), .A1(n126), .B0(n110), .B1(n78), .C0(n109), .C1(
        n108), .Y(n112) );
  OAI211XL U63 ( .A0(n107), .A1(n131), .B0(n2), .C0(addr[6]), .Y(n113) );
  OAI21XL U64 ( .A0(n1), .A1(addr[1]), .B0(n13), .Y(n81) );
  AOI221XL U65 ( .A0(n87), .A1(n78), .B0(n88), .B1(n126), .C0(n86), .Y(n90) );
  OAI211X1 U66 ( .A0(n85), .A1(n16), .B0(n84), .C0(n83), .Y(n86) );
  AOI222XL U67 ( .A0(n82), .A1(n78), .B0(n108), .B1(n107), .C0(n131), .C1(n79), 
        .Y(n85) );
  OAI21XL U68 ( .A0(n92), .A1(n7), .B0(addr[4]), .Y(n84) );
  AOI221XL U69 ( .A0(n126), .A1(n15), .B0(addr[3]), .B1(n127), .C0(n97), .Y(
        n98) );
  OAI22X1 U70 ( .A0(n5), .A1(n18), .B0(n20), .B1(n10), .Y(n97) );
  OAI211X1 U71 ( .A0(n14), .A1(n18), .B0(n119), .C0(n118), .Y(dout[3]) );
  AOI32XL U72 ( .A0(n126), .A1(n4), .A2(n103), .B0(n109), .B1(n110), .Y(n119)
         );
  AOI22XL U73 ( .A0(n117), .A1(n19), .B0(addr[5]), .B1(n116), .Y(n118) );
  AOI221XL U74 ( .A0(n122), .A1(n126), .B0(n96), .B1(n109), .C0(n8), .Y(n89)
         );
  AOI221XL U75 ( .A0(n131), .A1(n81), .B0(n95), .B1(n123), .C0(n80), .Y(n91)
         );
  NAND4X1 U76 ( .A(n102), .B(n114), .C(n101), .D(n100), .Y(dout[2]) );
  NAND3XL U77 ( .A(n3), .B(n125), .C(n103), .Y(n102) );
  AOI2BB2XL U78 ( .B0(addr[5]), .B1(n99), .A0N(addr[5]), .A1N(n98), .Y(n100)
         );
  OAI221X1 U79 ( .A0(n134), .A1(n19), .B0(n3), .B1(n133), .C0(n132), .Y(
        dout[4]) );
  AOI32XL U80 ( .A0(n131), .A1(n11), .A2(n1), .B0(n130), .B1(n19), .Y(n132) );
  AOI222XL U81 ( .A0(n15), .A1(n123), .B0(n122), .B1(addr[1]), .C0(n121), .C1(
        n6), .Y(n134) );
  CLKINVX3 U82 ( .A(n3), .Y(n76) );
  CLKINVX3 U83 ( .A(addr[3]), .Y(n78) );
endmodule


module sbox4_8 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126;

  OAI32X4 U12 ( .A0(n12), .A1(n2), .A2(addr[2]), .B0(n71), .B1(n108), .Y(n123)
         );
  OAI222X4 U20 ( .A0(addr[2]), .A1(n92), .B0(n106), .B1(n91), .C0(n90), .C1(
        n16), .Y(dout[2]) );
  OAI222X4 U33 ( .A0(addr[4]), .A1(n106), .B0(n72), .B1(n108), .C0(n2), .C1(
        n118), .Y(n83) );
  NAND2X2 U34 ( .A(addr[4]), .B(n2), .Y(n108) );
  NOR2X2 U43 ( .A(n14), .B(addr[4]), .Y(n113) );
  NOR2X2 U45 ( .A(n71), .B(n2), .Y(n111) );
  NAND2X2 U51 ( .A(n72), .B(n8), .Y(n118) );
  NOR2X2 U52 ( .A(n13), .B(addr[5]), .Y(n97) );
  NAND2X2 U53 ( .A(addr[6]), .B(addr[1]), .Y(n85) );
  NAND2X2 U54 ( .A(addr[1]), .B(n8), .Y(n116) );
  NOR2X2 U55 ( .A(n115), .B(n71), .Y(n121) );
  NAND2X2 U56 ( .A(n14), .B(n13), .Y(n115) );
  NAND2X2 U57 ( .A(addr[5]), .B(n13), .Y(n96) );
  NAND2X2 U58 ( .A(addr[6]), .B(n72), .Y(n106) );
  OAI222X1 U1 ( .A0(n12), .A1(n85), .B0(n97), .B1(n116), .C0(n13), .C1(n118), 
        .Y(n73) );
  CLKINVX1 U2 ( .A(n116), .Y(n7) );
  OAI31X4 U3 ( .A0(n118), .A1(n71), .A2(n13), .B0(n117), .Y(n119) );
  CLKINVX1 U4 ( .A(n14), .Y(n1) );
  CLKBUFX3 U5 ( .A(addr[3]), .Y(n2) );
  OAI221X1 U6 ( .A0(addr[2]), .A1(n80), .B0(n118), .B1(n105), .C0(n79), .Y(
        dout[1]) );
  INVX4 U7 ( .A(addr[5]), .Y(n71) );
  OAI31X1 U8 ( .A0(n108), .A1(addr[5]), .A2(n9), .B0(n107), .Y(n109) );
  AOI222XL U9 ( .A0(n13), .A1(n8), .B0(n113), .B1(n72), .C0(addr[1]), .C1(n14), 
        .Y(n114) );
  OAI222X1 U10 ( .A0(addr[1]), .A1(n84), .B0(n85), .B1(n74), .C0(n14), .C1(
        n107), .Y(n75) );
  NAND2XL U11 ( .A(n1), .B(addr[5]), .Y(n84) );
  AOI211XL U13 ( .A0(n83), .A1(n71), .B0(n82), .C0(n4), .Y(n92) );
  NAND2XL U14 ( .A(n13), .B(n71), .Y(n74) );
  CLKINVX1 U15 ( .A(n118), .Y(n3) );
  CLKINVX1 U16 ( .A(n115), .Y(n11) );
  CLKINVX1 U17 ( .A(n112), .Y(n6) );
  OAI21X1 U18 ( .A0(n7), .A1(n9), .B0(n16), .Y(n112) );
  AOI22X1 U19 ( .A0(n10), .A1(n111), .B0(n9), .B1(n113), .Y(n93) );
  OAI211X1 U21 ( .A0(n72), .A1(n115), .B0(n93), .C0(n5), .Y(n94) );
  CLKINVX1 U22 ( .A(n85), .Y(n10) );
  NAND2X1 U23 ( .A(n97), .B(n14), .Y(n105) );
  NAND2X1 U24 ( .A(n113), .B(n3), .Y(n98) );
  NAND2X1 U25 ( .A(n7), .B(n97), .Y(n107) );
  NAND2X1 U26 ( .A(n118), .B(n85), .Y(n110) );
  OAI21XL U27 ( .A0(n11), .A1(n71), .B0(n108), .Y(n95) );
  CLKINVX1 U28 ( .A(n84), .Y(n15) );
  CLKINVX1 U29 ( .A(addr[2]), .Y(n16) );
  OAI31X1 U30 ( .A0(n13), .A1(addr[6]), .A2(n71), .B0(n87), .Y(n88) );
  OAI21XL U31 ( .A0(n113), .A1(n12), .B0(n10), .Y(n87) );
  OAI211X1 U32 ( .A0(n76), .A1(n13), .B0(n98), .C0(n5), .Y(n77) );
  AOI222XL U35 ( .A0(addr[5]), .A1(addr[6]), .B0(n111), .B1(addr[1]), .C0(n9), 
        .C1(n2), .Y(n76) );
  NAND3XL U36 ( .A(n10), .B(n14), .C(addr[4]), .Y(n117) );
  OAI22XL U37 ( .A0(n116), .A1(n115), .B0(n1), .B1(n112), .Y(n78) );
  CLKINVX3 U38 ( .A(addr[4]), .Y(n13) );
  OAI2BB2XL U39 ( .B0(n115), .B1(n106), .A0N(n71), .A1N(n86), .Y(n89) );
  OAI221XL U40 ( .A0(n116), .A1(addr[4]), .B0(n108), .B1(addr[1]), .C0(n117), 
        .Y(n86) );
  CLKINVX1 U41 ( .A(addr[6]), .Y(n8) );
  CLKINVX1 U42 ( .A(n81), .Y(n4) );
  OAI21XL U44 ( .A0(n96), .A1(n118), .B0(n93), .Y(n82) );
  NAND3X1 U46 ( .A(n101), .B(n100), .C(n99), .Y(n102) );
  AOI32X1 U47 ( .A0(n96), .A1(n14), .A2(n7), .B0(n10), .B1(n95), .Y(n101) );
  AOI2BB2XL U48 ( .B0(n72), .B1(n121), .A0N(n98), .A1N(addr[5]), .Y(n99) );
  OAI21XL U49 ( .A0(n97), .A1(n12), .B0(n9), .Y(n100) );
  AOI2BB2XL U50 ( .B0(n9), .B1(n123), .A0N(n122), .A1N(n16), .Y(n124) );
  AOI211XL U59 ( .A0(n9), .A1(n121), .B0(n120), .C0(n119), .Y(n122) );
  OAI22XL U60 ( .A0(n116), .A1(n115), .B0(addr[5]), .B1(n114), .Y(n120) );
  CLKINVX1 U61 ( .A(n75), .Y(n5) );
  AOI32XL U62 ( .A0(n7), .A1(n96), .A2(n1), .B0(addr[1]), .B1(n121), .Y(n81)
         );
  AOI222XL U63 ( .A0(n9), .A1(n12), .B0(n121), .B1(n116), .C0(n2), .C1(n73), 
        .Y(n80) );
  AOI22XL U64 ( .A0(n78), .A1(n71), .B0(addr[2]), .B1(n77), .Y(n79) );
  NAND2XL U65 ( .A(n111), .B(addr[4]), .Y(n91) );
  AOI211X1 U66 ( .A0(n15), .A1(n110), .B0(n89), .C0(n88), .Y(n90) );
  OAI211X1 U67 ( .A0(n106), .A1(n105), .B0(n104), .C0(n103), .Y(dout[3]) );
  AOI32X1 U68 ( .A0(n2), .A1(n12), .A2(n7), .B0(n94), .B1(n16), .Y(n104) );
  AOI22XL U69 ( .A0(addr[2]), .A1(n102), .B0(n3), .B1(n123), .Y(n103) );
  OAI211X1 U70 ( .A0(addr[2]), .A1(n126), .B0(n125), .C0(n124), .Y(dout[4]) );
  AOI32X1 U71 ( .A0(n10), .A1(n12), .A2(n2), .B0(n6), .B1(n15), .Y(n125) );
  AOI221XL U72 ( .A0(n3), .A1(n111), .B0(n11), .B1(n110), .C0(n109), .Y(n126)
         );
  CLKINVX3 U73 ( .A(n106), .Y(n9) );
  CLKINVX3 U74 ( .A(n96), .Y(n12) );
  CLKINVX3 U75 ( .A(n2), .Y(n14) );
  CLKINVX3 U76 ( .A(addr[1]), .Y(n72) );
endmodule


module sbox5_8 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121;

  OAI222X4 U18 ( .A0(addr[3]), .A1(n106), .B0(n13), .B1(n90), .C0(n16), .C1(n8), .Y(n93) );
  OAI22X2 U40 ( .A0(addr[5]), .A1(n106), .B0(n14), .B1(n114), .Y(n116) );
  NOR2X2 U41 ( .A(n3), .B(addr[3]), .Y(n102) );
  NAND2X2 U45 ( .A(addr[6]), .B(n8), .Y(n114) );
  NAND2X2 U50 ( .A(n8), .B(n13), .Y(n110) );
  NAND2X2 U52 ( .A(addr[1]), .B(n13), .Y(n113) );
  NAND2X2 U54 ( .A(addr[1]), .B(addr[6]), .Y(n106) );
  NAND2X2 U55 ( .A(addr[3]), .B(n16), .Y(n121) );
  CLKINVX1 U1 ( .A(addr[5]), .Y(n1) );
  AOI221XL U2 ( .A0(n93), .A1(n1), .B0(n9), .B1(n68), .C0(n92), .Y(n105) );
  INVX3 U3 ( .A(addr[5]), .Y(n14) );
  OAI221X4 U4 ( .A0(n111), .A1(n110), .B0(n121), .B1(n114), .C0(n109), .Y(n112) );
  OAI221X4 U5 ( .A0(n16), .A1(n114), .B0(n14), .B1(n113), .C0(n120), .Y(n115)
         );
  OAI221X4 U6 ( .A0(n107), .A1(n121), .B0(n111), .B1(n113), .C0(n85), .Y(n86)
         );
  OAI31X1 U7 ( .A0(n70), .A1(addr[5]), .A2(addr[1]), .B0(n81), .Y(n73) );
  OAI32X1 U8 ( .A0(n114), .A1(addr[5]), .A2(n3), .B0(n15), .B1(n107), .Y(n79)
         );
  AOI32XL U9 ( .A0(n68), .A1(n98), .A2(n11), .B0(n2), .B1(n73), .Y(n77) );
  CLKBUFX3 U10 ( .A(addr[4]), .Y(n2) );
  CLKINVX1 U11 ( .A(n81), .Y(n4) );
  NAND2X1 U12 ( .A(n5), .B(n68), .Y(n81) );
  CLKINVX1 U13 ( .A(n110), .Y(n7) );
  CLKXOR2X2 U14 ( .A(n70), .B(n14), .Y(n94) );
  AOI2BB1X1 U15 ( .A0N(n16), .A1N(n1), .B0(n68), .Y(n111) );
  NOR2X1 U16 ( .A(n121), .B(n14), .Y(n91) );
  NOR2BX1 U17 ( .AN(n116), .B(n90), .Y(n83) );
  NAND2X1 U19 ( .A(n7), .B(n14), .Y(n120) );
  CLKINVX1 U20 ( .A(n113), .Y(n11) );
  NAND2X1 U21 ( .A(n11), .B(n14), .Y(n107) );
  CLKINVX1 U22 ( .A(n121), .Y(n15) );
  OAI31X1 U23 ( .A0(n12), .A1(n68), .A2(n113), .B0(n99), .Y(n72) );
  CLKINVX1 U24 ( .A(n106), .Y(n9) );
  OAI2BB2XL U25 ( .B0(n1), .B1(n113), .A0N(n98), .A1N(n5), .Y(n101) );
  CLKINVX1 U26 ( .A(n114), .Y(n5) );
  CLKINVX1 U27 ( .A(n90), .Y(n69) );
  CLKINVX1 U28 ( .A(addr[1]), .Y(n8) );
  CLKINVX1 U29 ( .A(addr[3]), .Y(n70) );
  CLKINVX1 U30 ( .A(addr[6]), .Y(n13) );
  AOI211X1 U31 ( .A0(n91), .A1(addr[1]), .B0(n80), .C0(n79), .Y(n89) );
  OAI2BB2XL U32 ( .B0(n111), .B1(n106), .A0N(n94), .A1N(n7), .Y(n80) );
  AOI211X1 U33 ( .A0(n102), .A1(n84), .B0(n83), .C0(n82), .Y(n85) );
  OAI21XL U34 ( .A0(n13), .A1(n1), .B0(n106), .Y(n84) );
  NOR3XL U35 ( .A(n94), .B(n3), .C(n110), .Y(n82) );
  AOI222XL U36 ( .A0(n9), .A1(n69), .B0(addr[5]), .B1(n108), .C0(n10), .C1(n16), .Y(n109) );
  CLKINVX1 U37 ( .A(n107), .Y(n10) );
  OAI21XL U38 ( .A0(addr[6]), .A1(addr[3]), .B0(n106), .Y(n108) );
  NAND2X1 U39 ( .A(addr[3]), .B(n3), .Y(n90) );
  NAND2X1 U42 ( .A(n2), .B(addr[5]), .Y(n98) );
  NAND2X1 U43 ( .A(n3), .B(n70), .Y(n97) );
  OAI21XL U44 ( .A0(addr[1]), .A1(n97), .B0(n96), .Y(n103) );
  AOI33XL U46 ( .A0(n3), .A1(n95), .A2(addr[5]), .B0(n94), .B1(n16), .B2(
        addr[1]), .Y(n96) );
  OAI21XL U47 ( .A0(n8), .A1(n70), .B0(n114), .Y(n95) );
  OAI21XL U48 ( .A0(addr[6]), .A1(n121), .B0(n99), .Y(n100) );
  NAND2X1 U49 ( .A(n71), .B(n7), .Y(n99) );
  XOR2X1 U51 ( .A(n12), .B(n3), .Y(n71) );
  AOI2BB2XL U53 ( .B0(n102), .B1(n116), .A0N(n2), .A1N(n75), .Y(n76) );
  AOI211X1 U56 ( .A0(n6), .A1(n3), .B0(n74), .C0(n83), .Y(n75) );
  AO22XL U57 ( .A0(n11), .A1(n15), .B0(addr[6]), .B1(n102), .Y(n74) );
  CLKINVX1 U58 ( .A(n120), .Y(n6) );
  CLKINVX1 U59 ( .A(n2), .Y(n12) );
  AO22XL U60 ( .A0(n11), .A1(n69), .B0(addr[6]), .B1(n91), .Y(n92) );
  AOI222XL U61 ( .A0(n116), .A1(n16), .B0(addr[3]), .B1(n115), .C0(n11), .C1(
        n68), .Y(n117) );
  OAI221X1 U62 ( .A0(n2), .A1(n105), .B0(n110), .B1(n121), .C0(n104), .Y(
        dout[3]) );
  AOI222XL U63 ( .A0(n2), .A1(n103), .B0(n102), .B1(n101), .C0(n100), .C1(n1), 
        .Y(n104) );
  OAI211X1 U64 ( .A0(n2), .A1(n89), .B0(n88), .C0(n87), .Y(dout[2]) );
  AOI33XL U65 ( .A0(n15), .A1(n98), .A2(n5), .B0(n3), .B1(n94), .B2(n7), .Y(
        n88) );
  AOI222XL U66 ( .A0(n4), .A1(n14), .B0(n2), .B1(n86), .C0(n91), .C1(n9), .Y(
        n87) );
  OAI211X1 U67 ( .A0(n78), .A1(n14), .B0(n77), .C0(n76), .Y(dout[1]) );
  AOI221XL U68 ( .A0(n15), .A1(addr[1]), .B0(n9), .B1(n68), .C0(n72), .Y(n78)
         );
  OAI211X1 U69 ( .A0(n121), .A1(n120), .B0(n119), .C0(n118), .Y(dout[4]) );
  AOI32XL U70 ( .A0(n68), .A1(n114), .A2(addr[5]), .B0(n2), .B1(n112), .Y(n119) );
  AOI2BB2X1 U71 ( .B0(n4), .B1(n14), .A0N(n2), .A1N(n117), .Y(n118) );
  BUFX4 U72 ( .A(addr[2]), .Y(n3) );
  CLKINVX3 U73 ( .A(n3), .Y(n16) );
  CLKINVX3 U74 ( .A(n97), .Y(n68) );
endmodule


module sbox6_8 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147;

  NAND2X2 U39 ( .A(n138), .B(addr[3]), .Y(n147) );
  NOR2X2 U47 ( .A(n15), .B(n10), .Y(n138) );
  NOR2X2 U50 ( .A(n85), .B(n4), .Y(n119) );
  NOR2X2 U58 ( .A(n83), .B(n85), .Y(n125) );
  NAND2X2 U61 ( .A(n97), .B(n103), .Y(n112) );
  NOR2X2 U62 ( .A(n17), .B(addr[1]), .Y(n103) );
  NOR2X2 U63 ( .A(n83), .B(addr[3]), .Y(n97) );
  NAND2X2 U64 ( .A(n117), .B(n131), .Y(n140) );
  NOR2X2 U65 ( .A(n5), .B(addr[3]), .Y(n131) );
  NOR2X2 U66 ( .A(n11), .B(addr[6]), .Y(n117) );
  NOR2X1 U1 ( .A(n15), .B(addr[3]), .Y(n102) );
  OAI222X1 U2 ( .A0(n91), .A1(n18), .B0(n2), .B1(n82), .C0(addr[5]), .C1(n84), 
        .Y(n92) );
  CLKINVX1 U3 ( .A(n83), .Y(n1) );
  INVX4 U4 ( .A(n4), .Y(n83) );
  CLKBUFX3 U5 ( .A(addr[4]), .Y(n4) );
  CLKINVX1 U6 ( .A(n15), .Y(n2) );
  BUFX4 U7 ( .A(addr[2]), .Y(n5) );
  CLKINVX1 U8 ( .A(addr[3]), .Y(n3) );
  OAI22X1 U9 ( .A0(n85), .A1(n17), .B0(addr[1]), .B1(n84), .Y(n142) );
  AOI211X1 U10 ( .A0(n18), .A1(n85), .B0(n131), .C0(n143), .Y(n121) );
  INVX3 U11 ( .A(addr[3]), .Y(n85) );
  OAI221X1 U12 ( .A0(n17), .A1(n81), .B0(n85), .B1(n8), .C0(n86), .Y(n90) );
  INVX3 U13 ( .A(n96), .Y(n8) );
  OAI221X4 U14 ( .A0(n123), .A1(n13), .B0(n10), .B1(n18), .C0(n7), .Y(n124) );
  NOR2X4 U15 ( .A(addr[1]), .B(addr[6]), .Y(n130) );
  NOR2X4 U16 ( .A(n5), .B(addr[5]), .Y(n143) );
  INVX1 U17 ( .A(n130), .Y(n14) );
  CLKINVX1 U18 ( .A(n125), .Y(n81) );
  NAND2X1 U19 ( .A(n14), .B(n8), .Y(n105) );
  INVXL U20 ( .A(n121), .Y(n16) );
  CLKINVX1 U21 ( .A(n138), .Y(n9) );
  CLKINVX1 U22 ( .A(n117), .Y(n10) );
  CLKINVX1 U23 ( .A(n119), .Y(n84) );
  NOR2X1 U24 ( .A(n8), .B(n123), .Y(n144) );
  NOR2X1 U25 ( .A(n11), .B(n17), .Y(n96) );
  CLKINVX1 U26 ( .A(n103), .Y(n13) );
  OAI211X1 U27 ( .A0(n14), .A1(n81), .B0(n104), .C0(n112), .Y(n108) );
  OAI21XL U28 ( .A0(n103), .A1(n117), .B0(n102), .Y(n104) );
  OAI21XL U29 ( .A0(n132), .A1(n17), .B0(n3), .Y(n86) );
  AOI21X1 U30 ( .A0(n83), .A1(n102), .B0(n125), .Y(n91) );
  OAI2BB2XL U31 ( .B0(n143), .B1(n14), .A0N(n143), .A1N(n117), .Y(n118) );
  CLKINVX1 U32 ( .A(n122), .Y(n7) );
  CLKINVX1 U33 ( .A(n126), .Y(n12) );
  CLKINVX1 U34 ( .A(n97), .Y(n82) );
  NAND2BX1 U35 ( .AN(n144), .B(n137), .Y(n107) );
  CLKINVX1 U36 ( .A(addr[1]), .Y(n11) );
  NOR2X1 U37 ( .A(n8), .B(n2), .Y(n122) );
  NOR2X1 U38 ( .A(addr[1]), .B(n1), .Y(n132) );
  OAI22X1 U40 ( .A0(n84), .A1(n10), .B0(n5), .B1(n12), .Y(n88) );
  NAND2X1 U41 ( .A(n5), .B(n18), .Y(n123) );
  NAND4X1 U42 ( .A(n147), .B(n140), .C(n100), .D(n99), .Y(n101) );
  AOI222XL U43 ( .A0(n98), .A1(n15), .B0(n102), .B1(n130), .C0(n97), .C1(n105), 
        .Y(n99) );
  NAND3X1 U44 ( .A(n5), .B(n84), .C(n96), .Y(n100) );
  OAI221X1 U45 ( .A0(n85), .A1(n13), .B0(n84), .B1(n17), .C0(n12), .Y(n98) );
  AOI22X1 U46 ( .A0(n4), .A1(n115), .B0(addr[5]), .B1(n114), .Y(n129) );
  OAI21XL U48 ( .A0(n121), .A1(n14), .B0(n147), .Y(n115) );
  OAI21XL U49 ( .A0(n113), .A1(n15), .B0(n112), .Y(n114) );
  AOI221XL U51 ( .A0(n119), .A1(n11), .B0(n130), .B1(addr[3]), .C0(n111), .Y(
        n113) );
  OAI22XL U52 ( .A0(n10), .A1(n83), .B0(addr[3]), .B1(n8), .Y(n111) );
  AOI211X1 U53 ( .A0(n4), .A1(n135), .B0(n134), .C0(n133), .Y(n136) );
  OA21XL U54 ( .A0(n3), .A1(n2), .B0(n132), .Y(n133) );
  OAI2BB2XL U55 ( .B0(n1), .B1(n7), .A0N(n131), .A1N(n130), .Y(n134) );
  OAI22X1 U56 ( .A0(n5), .A1(n10), .B0(n15), .B1(n8), .Y(n135) );
  CLKINVX3 U57 ( .A(addr[5]), .Y(n18) );
  AOI2BB2X1 U59 ( .B0(n5), .B1(n130), .A0N(n2), .A1N(n13), .Y(n137) );
  NOR2X1 U60 ( .A(n13), .B(n1), .Y(n126) );
  AOI2BB2XL U67 ( .B0(n143), .B1(n90), .A0N(n89), .A1N(n18), .Y(n94) );
  AOI211X1 U68 ( .A0(n122), .A1(n4), .B0(n88), .C0(n87), .Y(n89) );
  OAI32X1 U69 ( .A0(n13), .A1(n85), .A2(n15), .B0(n9), .B1(n82), .Y(n87) );
  NAND3X1 U70 ( .A(n147), .B(n140), .C(n139), .Y(n141) );
  AOI32X1 U71 ( .A0(n5), .A1(n11), .A2(n4), .B0(n138), .B1(n83), .Y(n139) );
  AO22XL U72 ( .A0(n143), .A1(n1), .B0(n116), .B1(n83), .Y(n120) );
  OAI21XL U73 ( .A0(n2), .A1(n18), .B0(n123), .Y(n116) );
  CLKINVX1 U74 ( .A(n106), .Y(n6) );
  AOI32XL U75 ( .A0(n105), .A1(n83), .A2(n3), .B0(addr[1]), .B1(n125), .Y(n106) );
  OAI211X1 U76 ( .A0(n83), .A1(n140), .B0(n110), .C0(n109), .Y(dout[2]) );
  AOI222XL U77 ( .A0(n108), .A1(n18), .B0(n143), .B1(n6), .C0(n119), .C1(n107), 
        .Y(n109) );
  AOI2BB2XL U78 ( .B0(addr[5]), .B1(n101), .A0N(n15), .A1N(n112), .Y(n110) );
  OAI211X1 U79 ( .A0(n1), .A1(n147), .B0(n146), .C0(n145), .Y(dout[4]) );
  AOI222XL U80 ( .A0(n144), .A1(n85), .B0(n143), .B1(n142), .C0(n141), .C1(n18), .Y(n145) );
  OA22X1 U81 ( .A0(n81), .A1(n137), .B0(n136), .B1(n18), .Y(n146) );
  NAND3X1 U82 ( .A(n129), .B(n128), .C(n127), .Y(dout[3]) );
  AOI32XL U83 ( .A0(n120), .A1(n85), .A2(addr[1]), .B0(n119), .B1(n118), .Y(
        n128) );
  AOI222XL U84 ( .A0(n144), .A1(n83), .B0(n126), .B1(n16), .C0(n125), .C1(n124), .Y(n127) );
  NAND3BX1 U85 ( .AN(n95), .B(n94), .C(n93), .Y(dout[1]) );
  OAI222X1 U86 ( .A0(n140), .A1(n4), .B0(n112), .B1(n15), .C0(n8), .C1(n91), 
        .Y(n95) );
  AOI32XL U87 ( .A0(addr[1]), .A1(n18), .A2(n125), .B0(n130), .B1(n92), .Y(n93) );
  CLKINVX3 U88 ( .A(n5), .Y(n15) );
  CLKINVX3 U89 ( .A(addr[6]), .Y(n17) );
endmodule


module sbox7_8 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148;

  OAI222X4 U19 ( .A0(n86), .A1(n129), .B0(n4), .B1(n18), .C0(addr[1]), .C1(n8), 
        .Y(n122) );
  OAI33X4 U33 ( .A0(addr[1]), .A1(n4), .A2(n5), .B0(n84), .B1(n6), .B2(n14), 
        .Y(n97) );
  NOR2X2 U44 ( .A(n17), .B(n4), .Y(n116) );
  NOR2X2 U48 ( .A(addr[1]), .B(addr[6]), .Y(n136) );
  NOR2X2 U51 ( .A(n20), .B(n17), .Y(n125) );
  NOR2X2 U52 ( .A(n84), .B(addr[3]), .Y(n131) );
  NOR2X2 U58 ( .A(n93), .B(n124), .Y(n142) );
  NOR2X2 U60 ( .A(n85), .B(addr[1]), .Y(n93) );
  NOR2X2 U62 ( .A(n12), .B(n3), .Y(n137) );
  NOR2X2 U65 ( .A(n85), .B(n87), .Y(n140) );
  NAND2X1 U1 ( .A(n3), .B(n4), .Y(n119) );
  CLKBUFX3 U2 ( .A(addr[4]), .Y(n4) );
  CLKINVX1 U3 ( .A(n12), .Y(n1) );
  CLKINVX1 U4 ( .A(n6), .Y(n2) );
  CLKBUFX3 U5 ( .A(addr[2]), .Y(n5) );
  OAI22X1 U6 ( .A0(addr[1]), .A1(n8), .B0(n5), .B1(n113), .Y(n100) );
  OAI31X1 U7 ( .A0(n17), .A1(n12), .A2(n87), .B0(n117), .Y(n121) );
  OAI22X1 U8 ( .A0(n4), .A1(n20), .B0(addr[3]), .B1(n11), .Y(n103) );
  NOR2X4 U9 ( .A(n87), .B(addr[6]), .Y(n124) );
  AOI211XL U10 ( .A0(n5), .A1(n83), .B0(n131), .C0(n130), .Y(n132) );
  NOR3XL U11 ( .A(n86), .B(addr[3]), .C(n2), .Y(n130) );
  OAI21XL U12 ( .A0(n3), .A1(n1), .B0(n119), .Y(n89) );
  BUFX4 U13 ( .A(addr[5]), .Y(n3) );
  AOI221XL U14 ( .A0(n140), .A1(n89), .B0(n109), .B1(n83), .C0(n88), .Y(n96)
         );
  CLKINVX1 U15 ( .A(n140), .Y(n84) );
  OAI2BB2XL U16 ( .B0(n142), .B1(n11), .A0N(n141), .A1N(n140), .Y(n143) );
  CLKINVX1 U17 ( .A(n125), .Y(n16) );
  CLKINVX1 U18 ( .A(n142), .Y(n83) );
  NAND2X1 U20 ( .A(n16), .B(n19), .Y(n105) );
  CLKINVX1 U21 ( .A(n123), .Y(n7) );
  CLKINVX1 U22 ( .A(n109), .Y(n10) );
  NAND2X1 U23 ( .A(n124), .B(n17), .Y(n113) );
  CLKINVX1 U24 ( .A(n137), .Y(n11) );
  NOR2X1 U25 ( .A(n11), .B(n17), .Y(n109) );
  CLKINVX1 U26 ( .A(n136), .Y(n86) );
  OAI22XL U27 ( .A0(n137), .A1(n18), .B0(n87), .B1(n10), .Y(n146) );
  OAI21X1 U28 ( .A0(n12), .A1(n16), .B0(n129), .Y(n141) );
  NAND2X1 U29 ( .A(n116), .B(n20), .Y(n129) );
  CLKINVX1 U30 ( .A(n93), .Y(n21) );
  OAI21XL U31 ( .A0(n119), .A1(n21), .B0(n118), .Y(n120) );
  OAI21XL U32 ( .A0(n125), .A1(n137), .B0(n124), .Y(n118) );
  NOR2X1 U34 ( .A(n20), .B(n8), .Y(n123) );
  CLKINVX1 U35 ( .A(n145), .Y(n8) );
  OAI22XL U36 ( .A0(n137), .A1(n113), .B0(n85), .B1(n7), .Y(n88) );
  CLKINVX1 U37 ( .A(n116), .Y(n14) );
  CLKINVX1 U38 ( .A(n131), .Y(n18) );
  CLKINVX1 U39 ( .A(n134), .Y(n19) );
  NOR2XL U40 ( .A(n125), .B(n12), .Y(n110) );
  CLKINVX1 U41 ( .A(n119), .Y(n13) );
  CLKINVX1 U42 ( .A(n103), .Y(n9) );
  OA21XL U43 ( .A0(n15), .A1(n21), .B0(n117), .Y(n102) );
  CLKINVX1 U45 ( .A(n105), .Y(n15) );
  OAI2BB1XL U46 ( .A0N(n103), .A1N(n124), .B0(n102), .Y(n104) );
  OAI22X1 U47 ( .A0(n20), .A1(n14), .B0(n4), .B1(n19), .Y(n112) );
  NOR4X1 U49 ( .A(n4), .B(addr[3]), .C(n87), .D(n6), .Y(n99) );
  XNOR2X1 U50 ( .A(addr[6]), .B(n5), .Y(n101) );
  AOI211X1 U53 ( .A0(n116), .A1(addr[6]), .B0(n115), .C0(n114), .Y(n128) );
  OAI222X1 U54 ( .A0(n111), .A1(n84), .B0(n110), .B1(n21), .C0(n86), .C1(n10), 
        .Y(n115) );
  OAI2BB2XL U55 ( .B0(n13), .B1(n113), .A0N(n87), .A1N(n112), .Y(n114) );
  OA21XL U56 ( .A0(n17), .A1(n3), .B0(n7), .Y(n111) );
  NAND2X1 U57 ( .A(n5), .B(n136), .Y(n133) );
  CLKINVX1 U59 ( .A(addr[6]), .Y(n85) );
  AOI211X1 U61 ( .A0(n131), .A1(n3), .B0(n92), .C0(n91), .Y(n95) );
  OAI221X1 U63 ( .A0(n87), .A1(n8), .B0(n84), .B1(n11), .C0(n102), .Y(n92) );
  OAI31X1 U64 ( .A0(n17), .A1(n12), .A2(n86), .B0(n90), .Y(n91) );
  AO21XL U66 ( .A0(n119), .A1(n129), .B0(addr[6]), .Y(n90) );
  NOR2X1 U67 ( .A(n12), .B(addr[3]), .Y(n145) );
  AOI21XL U68 ( .A0(addr[3]), .A1(n98), .B0(n97), .Y(n108) );
  OAI2BB1XL U69 ( .A0N(n6), .A1N(n124), .B0(n133), .Y(n98) );
  NAND3X1 U70 ( .A(n136), .B(n17), .C(n3), .Y(n117) );
  NOR2X1 U71 ( .A(addr[3]), .B(n3), .Y(n134) );
  OAI21X1 U72 ( .A0(n5), .A1(n142), .B0(n133), .Y(n138) );
  OAI22XL U73 ( .A0(n142), .A1(n14), .B0(n1), .B1(n132), .Y(n135) );
  AO21X1 U74 ( .A0(n139), .A1(n20), .B0(n138), .Y(n144) );
  OAI21XL U75 ( .A0(n2), .A1(n87), .B0(n21), .Y(n139) );
  OAI221X1 U76 ( .A0(n96), .A1(n6), .B0(n5), .B1(n95), .C0(n94), .Y(dout[1])
         );
  AOI2BB2X1 U77 ( .B0(n93), .B1(n112), .A0N(n133), .A1N(n9), .Y(n94) );
  OAI211X1 U78 ( .A0(n128), .A1(n6), .B0(n127), .C0(n126), .Y(dout[3]) );
  AOI32XL U79 ( .A0(n125), .A1(n1), .A2(n124), .B0(n123), .B1(n136), .Y(n126)
         );
  OAI31X1 U80 ( .A0(n122), .A1(n121), .A2(n120), .B0(n6), .Y(n127) );
  OAI221X1 U81 ( .A0(n3), .A1(n108), .B0(n107), .B1(n20), .C0(n106), .Y(
        dout[2]) );
  AOI32XL U82 ( .A0(n105), .A1(n6), .A2(n140), .B0(n2), .B1(n104), .Y(n106) );
  AOI211X1 U83 ( .A0(n101), .A1(n4), .B0(n100), .C0(n99), .Y(n107) );
  NAND2X1 U84 ( .A(n148), .B(n147), .Y(dout[4]) );
  AOI222XL U85 ( .A0(n136), .A1(n141), .B0(n3), .B1(n135), .C0(n134), .C1(n138), .Y(n148) );
  AOI222XL U86 ( .A0(n5), .A1(n146), .B0(n145), .B1(n144), .C0(n143), .C1(n6), 
        .Y(n147) );
  CLKINVX3 U87 ( .A(n5), .Y(n6) );
  CLKINVX3 U88 ( .A(n4), .Y(n12) );
  CLKINVX3 U89 ( .A(addr[3]), .Y(n17) );
  CLKINVX3 U90 ( .A(n3), .Y(n20) );
  CLKINVX3 U91 ( .A(addr[1]), .Y(n87) );
endmodule


module sbox8_8 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132;

  NAND2X2 U41 ( .A(addr[6]), .B(n15), .Y(n131) );
  NAND2X2 U48 ( .A(addr[4]), .B(n11), .Y(n123) );
  NAND2X2 U49 ( .A(n2), .B(n12), .Y(n87) );
  NAND2X2 U50 ( .A(addr[1]), .B(n75), .Y(n124) );
  NAND2X2 U54 ( .A(addr[2]), .B(n9), .Y(n116) );
  NAND2X2 U60 ( .A(addr[6]), .B(addr[1]), .Y(n105) );
  NAND2X2 U61 ( .A(n15), .B(n75), .Y(n108) );
  OAI32X1 U1 ( .A0(n75), .A1(addr[4]), .A2(n92), .B0(n115), .B1(n108), .Y(n96)
         );
  OAI31X1 U2 ( .A0(n123), .A1(addr[6]), .A2(n116), .B0(n109), .Y(n110) );
  OAI221X1 U3 ( .A0(n105), .A1(n87), .B0(addr[4]), .B1(n108), .C0(n86), .Y(n90) );
  NAND2X4 U4 ( .A(addr[4]), .B(n2), .Y(n115) );
  AOI222X1 U5 ( .A0(n88), .A1(addr[2]), .B0(n12), .B1(n4), .C0(n5), .C1(n92), 
        .Y(n114) );
  OAI222X1 U6 ( .A0(addr[2]), .A1(n126), .B0(n11), .B1(n125), .C0(n124), .C1(
        n123), .Y(n127) );
  AOI32XL U7 ( .A0(n74), .A1(n7), .A2(n2), .B0(n14), .B1(n117), .Y(n130) );
  OA21XL U8 ( .A0(n5), .A1(n9), .B0(n121), .Y(n78) );
  INVXL U9 ( .A(n119), .Y(n3) );
  INVX3 U10 ( .A(n2), .Y(n11) );
  BUFX4 U11 ( .A(addr[3]), .Y(n2) );
  CLKBUFX3 U12 ( .A(addr[5]), .Y(n1) );
  CLKINVX1 U13 ( .A(n108), .Y(n14) );
  CLKINVX1 U14 ( .A(n107), .Y(n6) );
  CLKINVX1 U15 ( .A(n93), .Y(n10) );
  NAND2X1 U16 ( .A(n11), .B(n12), .Y(n93) );
  NAND2X1 U17 ( .A(n5), .B(n9), .Y(n121) );
  OAI21XL U18 ( .A0(n115), .A1(n9), .B0(n107), .Y(n77) );
  OAI21X1 U19 ( .A0(n12), .A1(n9), .B0(n123), .Y(n88) );
  OAI31XL U20 ( .A0(n115), .A1(n15), .A2(n116), .B0(n118), .Y(n94) );
  CLKINVX1 U21 ( .A(n131), .Y(n13) );
  NAND2X1 U22 ( .A(n7), .B(n11), .Y(n107) );
  OAI22XL U23 ( .A0(n116), .A1(n123), .B0(n7), .B1(n115), .Y(n117) );
  OAI22XL U24 ( .A0(n123), .A1(n108), .B0(n131), .B1(n93), .Y(n95) );
  OAI2BB2XL U25 ( .B0(n115), .B1(n131), .A0N(n88), .A1N(n16), .Y(n89) );
  AOI211XL U26 ( .A0(n108), .A1(n105), .B0(n12), .C0(n121), .Y(n85) );
  CLKINVX1 U27 ( .A(n124), .Y(n74) );
  OAI22XL U28 ( .A0(n7), .A1(n123), .B0(n78), .B1(n87), .Y(n81) );
  NAND2BX2 U29 ( .AN(n78), .B(n11), .Y(n120) );
  NAND2XL U30 ( .A(n115), .B(n93), .Y(n104) );
  OAI2BB2XL U31 ( .B0(n106), .B1(n105), .A0N(n104), .A1N(n74), .Y(n111) );
  NOR2BXL U32 ( .AN(n123), .B(n103), .Y(n106) );
  NAND3X1 U33 ( .A(n104), .B(n15), .C(n7), .Y(n84) );
  AO21X1 U34 ( .A0(n7), .A1(n16), .B0(n101), .Y(n102) );
  OAI33X1 U35 ( .A0(n75), .A1(n11), .A2(n100), .B0(n5), .B1(n103), .B2(n124), 
        .Y(n101) );
  OA22XL U36 ( .A0(n107), .A1(n131), .B0(n120), .B1(n124), .Y(n98) );
  CLKINVX1 U37 ( .A(n125), .Y(n8) );
  OAI21XL U38 ( .A0(n74), .A1(n13), .B0(addr[4]), .Y(n86) );
  NAND2X1 U39 ( .A(n1), .B(n5), .Y(n100) );
  OAI221X1 U40 ( .A0(n124), .A1(n121), .B0(addr[1]), .B1(n120), .C0(n3), .Y(
        n128) );
  OAI31XL U42 ( .A0(n5), .A1(n15), .A2(n11), .B0(n118), .Y(n119) );
  NAND2X1 U43 ( .A(n16), .B(addr[2]), .Y(n125) );
  NAND4XL U44 ( .A(n13), .B(n1), .C(n2), .D(addr[2]), .Y(n109) );
  NAND3X1 U45 ( .A(n7), .B(n75), .C(n2), .Y(n118) );
  OAI21XL U46 ( .A0(n1), .A1(n87), .B0(n114), .Y(n76) );
  OAI22XL U47 ( .A0(n108), .A1(n120), .B0(n79), .B1(n100), .Y(n80) );
  AOI221XL U51 ( .A0(n13), .A1(n11), .B0(n16), .B1(n2), .C0(n91), .Y(n79) );
  NOR2X1 U52 ( .A(n1), .B(n2), .Y(n103) );
  NOR2X1 U53 ( .A(n87), .B(addr[6]), .Y(n91) );
  NOR2X1 U55 ( .A(n11), .B(n1), .Y(n92) );
  CLKINVX1 U56 ( .A(n100), .Y(n4) );
  OA21XL U57 ( .A0(n1), .A1(n115), .B0(n120), .Y(n132) );
  AOI221XL U58 ( .A0(n14), .A1(n2), .B0(n16), .B1(addr[4]), .C0(n122), .Y(n126) );
  OAI22XL U59 ( .A0(n2), .A1(n15), .B0(addr[4]), .B1(n131), .Y(n122) );
  OAI211X1 U62 ( .A0(addr[2]), .A1(n99), .B0(n98), .C0(n97), .Y(dout[2]) );
  AOI221XL U63 ( .A0(addr[2]), .A1(n96), .B0(n1), .B1(n95), .C0(n94), .Y(n97)
         );
  AOI221XL U64 ( .A0(n91), .A1(n1), .B0(n90), .B1(n9), .C0(n89), .Y(n99) );
  OAI211X1 U65 ( .A0(n132), .A1(n131), .B0(n130), .C0(n129), .Y(dout[4]) );
  AOI222XL U66 ( .A0(n128), .A1(n12), .B0(n1), .B1(n127), .C0(n6), .C1(n16), 
        .Y(n129) );
  OAI211X1 U67 ( .A0(addr[1]), .A1(n114), .B0(n113), .C0(n112), .Y(dout[3]) );
  AOI221XL U68 ( .A0(n111), .A1(n5), .B0(n6), .B1(n14), .C0(n110), .Y(n112) );
  AOI2BB2XL U69 ( .B0(n102), .B1(n12), .A0N(n115), .A1N(n125), .Y(n113) );
  NAND4BX1 U70 ( .AN(n85), .B(n84), .C(n83), .D(n82), .Y(dout[1]) );
  AOI221XL U71 ( .A0(n13), .A1(n81), .B0(n10), .B1(n8), .C0(n80), .Y(n82) );
  AOI22X1 U72 ( .A0(n16), .A1(n77), .B0(n74), .B1(n76), .Y(n83) );
  CLKINVX3 U73 ( .A(addr[2]), .Y(n5) );
  CLKINVX3 U74 ( .A(n116), .Y(n7) );
  CLKINVX3 U75 ( .A(n1), .Y(n9) );
  CLKINVX3 U76 ( .A(addr[4]), .Y(n12) );
  CLKINVX3 U77 ( .A(addr[1]), .Y(n15) );
  CLKINVX3 U78 ( .A(n105), .Y(n16) );
  CLKINVX3 U79 ( .A(addr[6]), .Y(n75) );
endmodule


module crp_8 ( P, R, K_sub );
  output [1:32] P;
  input [1:32] R;
  input [1:48] K_sub;
  wire   n1;
  wire   [1:48] X;

  sbox1_8 u0 ( .addr(X[1:6]), .dout({P[9], P[17], P[23], P[31]}) );
  sbox2_8 u1 ( .addr({X[7], n1, X[9:12]}), .dout({P[13], P[28], P[2], P[18]})
         );
  sbox3_8 u2 ( .addr(X[13:18]), .dout({P[24], P[16], P[30], P[6]}) );
  sbox4_8 u3 ( .addr(X[19:24]), .dout({P[26], P[20], P[10], P[1]}) );
  sbox5_8 u4 ( .addr(X[25:30]), .dout({P[8], P[14], P[25], P[3]}) );
  sbox6_8 u5 ( .addr(X[31:36]), .dout({P[4], P[29], P[11], P[19]}) );
  sbox7_8 u6 ( .addr(X[37:42]), .dout({P[32], P[12], P[22], P[7]}) );
  sbox8_8 u7 ( .addr(X[43:48]), .dout({P[5], P[27], P[15], P[21]}) );
  XOR2X1 U1 ( .A(R[1]), .B(K_sub[2]), .Y(X[2]) );
  CLKXOR2X4 U2 ( .A(R[5]), .B(K_sub[6]), .Y(X[6]) );
  CLKXOR2X4 U3 ( .A(R[16]), .B(K_sub[25]), .Y(X[25]) );
  CLKXOR2X4 U4 ( .A(R[29]), .B(K_sub[42]), .Y(X[42]) );
  CLKXOR2X4 U5 ( .A(R[8]), .B(K_sub[11]), .Y(X[11]) );
  CLKXOR2X4 U6 ( .A(R[22]), .B(K_sub[33]), .Y(X[33]) );
  CLKXOR2X4 U7 ( .A(R[16]), .B(K_sub[23]), .Y(X[23]) );
  CLKXOR2X4 U8 ( .A(R[26]), .B(K_sub[39]), .Y(X[39]) );
  CLKXOR2X4 U9 ( .A(R[10]), .B(K_sub[15]), .Y(X[15]) );
  XNOR2X1 U10 ( .A(R[5]), .B(K_sub[8]), .Y(X[8]) );
  INVX3 U11 ( .A(X[8]), .Y(n1) );
  CLKXOR2X4 U12 ( .A(R[20]), .B(K_sub[31]), .Y(X[31]) );
  CLKXOR2X4 U13 ( .A(R[31]), .B(K_sub[46]), .Y(X[46]) );
  CLKXOR2X4 U14 ( .A(R[29]), .B(K_sub[44]), .Y(X[44]) );
  CLKXOR2X4 U15 ( .A(R[12]), .B(K_sub[19]), .Y(X[19]) );
  CLKXOR2X4 U16 ( .A(R[20]), .B(K_sub[29]), .Y(X[29]) );
  CLKXOR2X2 U17 ( .A(R[4]), .B(K_sub[5]), .Y(X[5]) );
  CLKXOR2X2 U18 ( .A(R[15]), .B(K_sub[22]), .Y(X[22]) );
  CLKXOR2X2 U19 ( .A(R[24]), .B(K_sub[35]), .Y(X[35]) );
  CLKXOR2X2 U20 ( .A(R[21]), .B(K_sub[30]), .Y(X[30]) );
  CLKXOR2X2 U21 ( .A(R[12]), .B(K_sub[17]), .Y(X[17]) );
  CLKXOR2X2 U22 ( .A(R[32]), .B(K_sub[1]), .Y(X[1]) );
  CLKXOR2X2 U23 ( .A(R[13]), .B(K_sub[20]), .Y(X[20]) );
  CLKXOR2X2 U24 ( .A(R[18]), .B(K_sub[27]), .Y(X[27]) );
  CLKXOR2X2 U25 ( .A(R[8]), .B(K_sub[13]), .Y(X[13]) );
  CLKXOR2X2 U26 ( .A(R[4]), .B(K_sub[7]), .Y(X[7]) );
  CLKXOR2X2 U27 ( .A(R[24]), .B(K_sub[37]), .Y(X[37]) );
  CLKXOR2X2 U28 ( .A(R[28]), .B(K_sub[43]), .Y(X[43]) );
  CLKXOR2X2 U29 ( .A(R[1]), .B(K_sub[48]), .Y(X[48]) );
  CLKXOR2X2 U30 ( .A(R[17]), .B(K_sub[24]), .Y(X[24]) );
  CLKXOR2X2 U31 ( .A(R[9]), .B(K_sub[12]), .Y(X[12]) );
  CLKXOR2X2 U32 ( .A(R[13]), .B(K_sub[18]), .Y(X[18]) );
  CLKXOR2X2 U33 ( .A(R[25]), .B(K_sub[36]), .Y(X[36]) );
  XOR2X1 U34 ( .A(R[23]), .B(K_sub[34]), .Y(X[34]) );
  XOR2X1 U35 ( .A(R[9]), .B(K_sub[14]), .Y(X[14]) );
  XOR2X1 U36 ( .A(R[30]), .B(K_sub[45]), .Y(X[45]) );
  XOR2X1 U37 ( .A(R[21]), .B(K_sub[32]), .Y(X[32]) );
  XOR2X1 U38 ( .A(R[25]), .B(K_sub[38]), .Y(X[38]) );
  XOR2X1 U39 ( .A(R[27]), .B(K_sub[40]), .Y(X[40]) );
  XOR2X1 U40 ( .A(R[3]), .B(K_sub[4]), .Y(X[4]) );
  XOR2X1 U41 ( .A(R[11]), .B(K_sub[16]), .Y(X[16]) );
  XOR2X1 U42 ( .A(R[7]), .B(K_sub[10]), .Y(X[10]) );
  XOR2X1 U43 ( .A(R[14]), .B(K_sub[21]), .Y(X[21]) );
  XOR2X1 U44 ( .A(R[6]), .B(K_sub[9]), .Y(X[9]) );
  XOR2X1 U45 ( .A(R[2]), .B(K_sub[3]), .Y(X[3]) );
  XOR2X1 U46 ( .A(R[28]), .B(K_sub[41]), .Y(X[41]) );
  XOR2X1 U47 ( .A(R[17]), .B(K_sub[26]), .Y(X[26]) );
  XOR2X1 U48 ( .A(R[32]), .B(K_sub[47]), .Y(X[47]) );
  XOR2X1 U49 ( .A(R[19]), .B(K_sub[28]), .Y(X[28]) );
endmodule


module sbox1_7 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127;

  OAI222X4 U13 ( .A0(addr[5]), .A1(n101), .B0(n1), .B1(n100), .C0(n99), .C1(
        n10), .Y(dout[3]) );
  OAI21X2 U42 ( .A0(n4), .A1(n112), .B0(n106), .Y(n123) );
  NAND2X2 U44 ( .A(addr[6]), .B(n72), .Y(n115) );
  NAND2X2 U48 ( .A(addr[1]), .B(n13), .Y(n114) );
  OAI22X2 U49 ( .A0(n6), .A1(n71), .B0(addr[5]), .B1(n120), .Y(n85) );
  NAND2X2 U50 ( .A(n3), .B(n6), .Y(n120) );
  NOR2X2 U51 ( .A(n6), .B(n3), .Y(n124) );
  NOR3X2 U55 ( .A(n2), .B(addr[6]), .C(n10), .Y(n102) );
  NOR2X2 U56 ( .A(n109), .B(n3), .Y(n93) );
  NAND2X2 U57 ( .A(addr[1]), .B(addr[6]), .Y(n109) );
  NAND2X2 U59 ( .A(n72), .B(n13), .Y(n112) );
  NOR2X1 U1 ( .A(n114), .B(n120), .Y(n104) );
  BUFX4 U2 ( .A(addr[4]), .Y(n2) );
  CLKBUFX3 U3 ( .A(addr[2]), .Y(n1) );
  OAI32X1 U4 ( .A0(n112), .A1(n2), .A2(n4), .B0(n115), .B1(n113), .Y(n80) );
  NOR2BXL U5 ( .AN(n118), .B(n1), .Y(n122) );
  CLKBUFX3 U6 ( .A(addr[2]), .Y(n4) );
  INVX3 U7 ( .A(addr[6]), .Y(n13) );
  OAI221X4 U8 ( .A0(n88), .A1(n71), .B0(addr[5]), .B1(n87), .C0(n86), .Y(
        dout[2]) );
  OAI221X4 U9 ( .A0(addr[5]), .A1(n127), .B0(n126), .B1(n71), .C0(n125), .Y(
        dout[4]) );
  OA21XL U10 ( .A0(n95), .A1(n115), .B0(n107), .Y(n119) );
  AOI222XL U11 ( .A0(n12), .A1(n1), .B0(n2), .B1(n110), .C0(n69), .C1(n10), 
        .Y(n111) );
  AOI2BB2X1 U12 ( .B0(n2), .B1(n69), .A0N(addr[4]), .A1N(n115), .Y(n91) );
  BUFX4 U14 ( .A(addr[3]), .Y(n3) );
  CLKINVX1 U15 ( .A(n112), .Y(n12) );
  CLKINVX1 U16 ( .A(n113), .Y(n7) );
  NAND2BX1 U17 ( .AN(n104), .B(n119), .Y(n84) );
  CLKXOR2X2 U18 ( .A(n8), .B(n10), .Y(n90) );
  NOR2X1 U19 ( .A(n6), .B(n8), .Y(n118) );
  OAI21XL U20 ( .A0(n8), .A1(n114), .B0(n91), .Y(n92) );
  NAND2X1 U21 ( .A(n93), .B(n6), .Y(n107) );
  NAND2X1 U22 ( .A(n10), .B(n8), .Y(n113) );
  OAI211X1 U23 ( .A0(n6), .A1(n114), .B0(n108), .C0(n107), .Y(n89) );
  CLKINVX1 U24 ( .A(n109), .Y(n69) );
  NAND2X1 U25 ( .A(n124), .B(n70), .Y(n108) );
  CLKINVX1 U26 ( .A(n114), .Y(n11) );
  CLKINVX1 U27 ( .A(n115), .Y(n70) );
  CLKINVX1 U28 ( .A(n95), .Y(n9) );
  AO22X1 U29 ( .A0(n90), .A1(n70), .B0(n8), .B1(n123), .Y(n76) );
  OAI31X1 U30 ( .A0(n10), .A1(n3), .A2(n72), .B0(n103), .Y(n105) );
  AOI31XL U31 ( .A0(n72), .A1(n10), .A2(n2), .B0(n102), .Y(n103) );
  AOI211X1 U32 ( .A0(n5), .A1(n4), .B0(n117), .C0(n116), .Y(n126) );
  CLKINVX1 U33 ( .A(n108), .Y(n5) );
  AOI211X1 U34 ( .A0(n115), .A1(n114), .B0(n113), .C0(n2), .Y(n116) );
  OAI22X1 U35 ( .A0(n120), .A1(n112), .B0(n111), .B1(n8), .Y(n117) );
  AOI211X1 U36 ( .A0(n69), .A1(n118), .B0(n81), .C0(n80), .Y(n88) );
  OAI22X1 U37 ( .A0(n91), .A1(n10), .B0(n3), .B1(n106), .Y(n81) );
  CLKINVX3 U38 ( .A(addr[5]), .Y(n71) );
  NAND2X1 U39 ( .A(n3), .B(n71), .Y(n95) );
  NAND2X1 U40 ( .A(n11), .B(n1), .Y(n106) );
  XOR2X1 U41 ( .A(n82), .B(n2), .Y(n83) );
  NAND2X1 U43 ( .A(n1), .B(n3), .Y(n82) );
  OAI22XL U45 ( .A0(n3), .A1(n72), .B0(n8), .B1(n112), .Y(n94) );
  AOI211XL U46 ( .A0(n98), .A1(n8), .B0(n97), .C0(n104), .Y(n99) );
  OAI22XL U47 ( .A0(n96), .A1(n6), .B0(n95), .B1(n109), .Y(n97) );
  OAI22XL U52 ( .A0(n13), .A1(n71), .B0(n2), .B1(addr[1]), .Y(n98) );
  AOI221XL U53 ( .A0(n9), .A1(addr[6]), .B0(addr[5]), .B1(n94), .C0(n93), .Y(
        n96) );
  OAI21XL U54 ( .A0(addr[1]), .A1(n120), .B0(n119), .Y(n121) );
  AOI221XL U58 ( .A0(n12), .A1(n118), .B0(n93), .B1(n71), .C0(n75), .Y(n78) );
  OAI31X1 U60 ( .A0(n71), .A1(n2), .A2(n74), .B0(n73), .Y(n75) );
  OA21XL U61 ( .A0(n3), .A1(n13), .B0(n109), .Y(n74) );
  OAI21XL U62 ( .A0(n124), .A1(n85), .B0(n11), .Y(n73) );
  OAI21XL U63 ( .A0(n1), .A1(n72), .B0(n109), .Y(n110) );
  INVX4 U64 ( .A(n4), .Y(n10) );
  AOI222XL U65 ( .A0(n124), .A1(n123), .B0(n122), .B1(addr[6]), .C0(n1), .C1(
        n121), .Y(n125) );
  NOR4BBX1 U66 ( .AN(n107), .BN(n106), .C(n105), .D(n104), .Y(n127) );
  AOI222XL U67 ( .A0(n12), .A1(n90), .B0(n89), .B1(n10), .C0(n123), .C1(n6), 
        .Y(n101) );
  AOI2BB2XL U68 ( .B0(addr[5]), .B1(n92), .A0N(n120), .A1N(addr[1]), .Y(n100)
         );
  AOI32X1 U69 ( .A0(n4), .A1(n85), .A2(n12), .B0(n84), .B1(n10), .Y(n86) );
  AOI222XL U70 ( .A0(n124), .A1(n72), .B0(n83), .B1(addr[1]), .C0(n7), .C1(n13), .Y(n87) );
  OAI221X1 U71 ( .A0(n79), .A1(n71), .B0(n4), .B1(n78), .C0(n77), .Y(dout[1])
         );
  AOI32XL U72 ( .A0(addr[6]), .A1(n85), .A2(n1), .B0(n76), .B1(n71), .Y(n77)
         );
  AOI221X1 U73 ( .A0(n12), .A1(n90), .B0(n4), .B1(n93), .C0(n102), .Y(n79) );
  CLKINVX3 U74 ( .A(n2), .Y(n6) );
  CLKINVX3 U75 ( .A(n3), .Y(n8) );
  CLKINVX3 U76 ( .A(addr[1]), .Y(n72) );
endmodule


module sbox2_7 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147;

  NAND2X2 U55 ( .A(n2), .B(n81), .Y(n136) );
  NAND2X2 U57 ( .A(addr[2]), .B(n15), .Y(n104) );
  NAND2X2 U60 ( .A(addr[5]), .B(addr[2]), .Y(n132) );
  NOR2X2 U61 ( .A(n7), .B(n4), .Y(n101) );
  NAND2X2 U62 ( .A(n6), .B(n13), .Y(n146) );
  NAND2X2 U63 ( .A(n3), .B(n83), .Y(n124) );
  NAND2X2 U64 ( .A(addr[6]), .B(n6), .Y(n122) );
  NAND2X2 U67 ( .A(n3), .B(n2), .Y(n133) );
  AOI222XL U1 ( .A0(n9), .A1(n8), .B0(n88), .B1(n83), .C0(n140), .C1(n4), .Y(
        n89) );
  CLKINVX1 U2 ( .A(n121), .Y(n7) );
  NOR2X1 U3 ( .A(n104), .B(n2), .Y(n141) );
  NOR2X1 U4 ( .A(n124), .B(n2), .Y(n140) );
  CLKBUFX4 U5 ( .A(addr[4]), .Y(n2) );
  CLKINVX1 U6 ( .A(addr[5]), .Y(n1) );
  INVX3 U7 ( .A(addr[5]), .Y(n15) );
  OAI211X4 U8 ( .A0(n147), .A1(n146), .B0(n145), .C0(n144), .Y(dout[4]) );
  NAND3XL U9 ( .A(n98), .B(n97), .C(n96), .Y(dout[1]) );
  NAND2X1 U10 ( .A(addr[1]), .B(addr[6]), .Y(n121) );
  CLKINVX2 U11 ( .A(addr[1]), .Y(n6) );
  OAI221X1 U12 ( .A0(addr[1]), .A1(n136), .B0(n133), .B1(n6), .C0(n87), .Y(n95) );
  NAND2X4 U13 ( .A(addr[1]), .B(n13), .Y(n114) );
  INVX3 U14 ( .A(addr[6]), .Y(n13) );
  NAND2XL U15 ( .A(n102), .B(n81), .Y(n109) );
  AOI211XL U16 ( .A0(n16), .A1(n95), .B0(n94), .C0(n93), .Y(n96) );
  AOI2BB2X1 U17 ( .B0(n15), .B1(n82), .A0N(n104), .A1N(n136), .Y(n117) );
  NOR3BXL U18 ( .AN(n135), .B(n134), .C(n9), .Y(n147) );
  BUFX4 U19 ( .A(addr[3]), .Y(n3) );
  NAND2X1 U20 ( .A(n9), .B(n7), .Y(n113) );
  CLKINVX1 U21 ( .A(n146), .Y(n4) );
  CLKINVX1 U22 ( .A(n115), .Y(n9) );
  CLKINVX1 U23 ( .A(n122), .Y(n5) );
  OAI31X1 U24 ( .A0(n124), .A1(n13), .A2(n15), .B0(n123), .Y(n128) );
  OAI21XL U25 ( .A0(n15), .A1(n6), .B0(n140), .Y(n123) );
  OAI22X1 U26 ( .A0(n122), .A1(n124), .B0(n101), .B1(n132), .Y(n84) );
  INVX1 U27 ( .A(n114), .Y(n8) );
  OAI22X1 U28 ( .A0(n122), .A1(n81), .B0(n10), .B1(n121), .Y(n129) );
  NAND3X1 U29 ( .A(n10), .B(n15), .C(n6), .Y(n111) );
  NAND2X1 U30 ( .A(n81), .B(n10), .Y(n115) );
  OAI21XL U31 ( .A0(n83), .A1(n133), .B0(n135), .Y(n85) );
  OAI22XL U32 ( .A0(n117), .A1(n146), .B0(n116), .B1(n132), .Y(n118) );
  AOI222XL U33 ( .A0(n8), .A1(n115), .B0(n11), .B1(n13), .C0(n9), .C1(n4), .Y(
        n116) );
  CLKINVX1 U34 ( .A(n104), .Y(n14) );
  OAI2BB2XL U35 ( .B0(n114), .B1(n135), .A0N(n126), .A1N(n11), .Y(n106) );
  OAI21XL U36 ( .A0(n112), .A1(n114), .B0(n111), .Y(n120) );
  OAI21XL U37 ( .A0(n133), .A1(n114), .B0(n113), .Y(n119) );
  CLKINVX1 U38 ( .A(n124), .Y(n82) );
  CLKINVX1 U39 ( .A(n136), .Y(n12) );
  CLKINVX1 U40 ( .A(n133), .Y(n11) );
  CLKINVX1 U41 ( .A(n132), .Y(n16) );
  AOI2BB1X1 U42 ( .A0N(n126), .A1N(n125), .B0(n136), .Y(n127) );
  OAI22XL U43 ( .A0(n104), .A1(n114), .B0(n101), .B1(n132), .Y(n102) );
  AO21XL U44 ( .A0(n83), .A1(n12), .B0(n141), .Y(n86) );
  AO21X1 U45 ( .A0(n81), .A1(n14), .B0(n140), .Y(n142) );
  NAND3X1 U46 ( .A(n83), .B(n10), .C(addr[5]), .Y(n135) );
  OAI22X1 U47 ( .A0(addr[5]), .A1(n121), .B0(n122), .B1(n15), .Y(n126) );
  AOI2BB1X1 U48 ( .A0N(n3), .A1N(n1), .B0(n12), .Y(n112) );
  NOR3X1 U49 ( .A(addr[1]), .B(addr[2]), .C(n15), .Y(n125) );
  AOI2BB1XL U50 ( .A0N(n92), .A1N(n91), .B0(addr[5]), .Y(n93) );
  OAI22XL U51 ( .A0(n117), .A1(n114), .B0(n89), .B1(n1), .Y(n94) );
  OAI31XL U52 ( .A0(n114), .A1(n2), .A2(n81), .B0(n90), .Y(n91) );
  OAI21XL U53 ( .A0(n11), .A1(n82), .B0(n5), .Y(n90) );
  NAND2X1 U54 ( .A(n8), .B(n2), .Y(n137) );
  OAI31XL U56 ( .A0(n101), .A1(n3), .A2(addr[2]), .B0(n113), .Y(n92) );
  OAI211X1 U58 ( .A0(n139), .A1(n15), .B0(n138), .C0(n137), .Y(n143) );
  NAND3X1 U59 ( .A(n10), .B(n15), .C(addr[6]), .Y(n138) );
  AOI2BB2X1 U65 ( .B0(n5), .B1(n81), .A0N(n6), .A1N(n136), .Y(n139) );
  OAI22XL U66 ( .A0(addr[5]), .A1(n133), .B0(n3), .B1(n132), .Y(n134) );
  OAI2BB2XL U68 ( .B0(n112), .B1(n122), .A0N(n1), .A1N(n99), .Y(n100) );
  OAI211X1 U69 ( .A0(n146), .A1(n2), .B0(n137), .C0(n113), .Y(n99) );
  NAND3X1 U70 ( .A(n5), .B(n10), .C(n3), .Y(n87) );
  AOI2BB2XL U71 ( .B0(n3), .B1(n105), .A0N(n137), .A1N(n132), .Y(n108) );
  OAI211XL U72 ( .A0(n104), .A1(n146), .B0(n103), .C0(n111), .Y(n105) );
  NAND3XL U73 ( .A(addr[5]), .B(n10), .C(n7), .Y(n103) );
  OAI22XL U74 ( .A0(n3), .A1(n114), .B0(n13), .B1(n115), .Y(n88) );
  NAND4X1 U75 ( .A(n110), .B(n109), .C(n108), .D(n107), .Y(dout[2]) );
  AOI32XL U76 ( .A0(addr[1]), .A1(addr[2]), .A2(n12), .B0(n100), .B1(n83), .Y(
        n110) );
  AOI221XL U77 ( .A0(n125), .A1(addr[4]), .B0(n141), .B1(n5), .C0(n106), .Y(
        n107) );
  AOI33XL U78 ( .A0(n5), .A1(n14), .A2(n2), .B0(n16), .B1(n146), .B2(n3), .Y(
        n145) );
  AOI222XL U79 ( .A0(n143), .A1(n83), .B0(n7), .B1(n142), .C0(n8), .C1(n141), 
        .Y(n144) );
  AOI32XL U80 ( .A0(n14), .A1(n6), .A2(n9), .B0(n4), .B1(n86), .Y(n97) );
  AOI22X1 U81 ( .A0(n7), .A1(n85), .B0(n2), .B1(n84), .Y(n98) );
  NAND2X1 U82 ( .A(n131), .B(n130), .Y(dout[3]) );
  AOI221XL U83 ( .A0(n120), .A1(n83), .B0(addr[2]), .B1(n119), .C0(n118), .Y(
        n131) );
  AOI211X1 U84 ( .A0(n14), .A1(n129), .B0(n128), .C0(n127), .Y(n130) );
  CLKINVX3 U85 ( .A(n2), .Y(n10) );
  CLKINVX3 U86 ( .A(n3), .Y(n81) );
  CLKINVX3 U87 ( .A(addr[2]), .Y(n83) );
endmodule


module sbox3_7 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133;

  NOR2X2 U35 ( .A(n13), .B(addr[3]), .Y(n108) );
  NOR2X2 U50 ( .A(addr[1]), .B(addr[6]), .Y(n107) );
  NOR2X2 U52 ( .A(n15), .B(n2), .Y(n87) );
  NOR2X2 U56 ( .A(n15), .B(n7), .Y(n94) );
  NOR2X1 U1 ( .A(n13), .B(n15), .Y(n106) );
  OAI221X1 U2 ( .A0(n124), .A1(n13), .B0(n3), .B1(addr[1]), .C0(n76), .Y(n104)
         );
  OAI22XL U3 ( .A0(n2), .A1(n7), .B0(n3), .B1(n11), .Y(n123) );
  BUFX4 U4 ( .A(addr[4]), .Y(n2) );
  CLKBUFX3 U5 ( .A(n7), .Y(n1) );
  OAI33X1 U6 ( .A0(n14), .A1(n125), .A2(n7), .B0(n13), .B1(n94), .B2(n119), 
        .Y(n79) );
  INVX3 U7 ( .A(n3), .Y(n7) );
  NOR2X1 U8 ( .A(n20), .B(n3), .Y(n91) );
  NOR2X1 U9 ( .A(n14), .B(n3), .Y(n121) );
  NOR2X1 U10 ( .A(n76), .B(n3), .Y(n95) );
  NOR2X1 U11 ( .A(n3), .B(n2), .Y(n110) );
  CLKBUFX4 U12 ( .A(addr[2]), .Y(n3) );
  OAI221X1 U13 ( .A0(addr[5]), .A1(n90), .B0(n89), .B1(n77), .C0(n88), .Y(
        dout[1]) );
  NOR2X4 U14 ( .A(n78), .B(n19), .Y(n124) );
  NOR2X4 U15 ( .A(addr[3]), .B(n2), .Y(n130) );
  NOR2X4 U16 ( .A(n19), .B(addr[6]), .Y(n125) );
  INVX3 U17 ( .A(addr[1]), .Y(n19) );
  NAND2XL U18 ( .A(n94), .B(n124), .Y(n132) );
  OAI211XL U19 ( .A0(n2), .A1(n8), .B0(n128), .C0(n127), .Y(n129) );
  NAND4XL U20 ( .A(n114), .B(n113), .C(n112), .D(n111), .Y(n115) );
  CLKINVX1 U21 ( .A(n132), .Y(n6) );
  INVX1 U22 ( .A(n124), .Y(n16) );
  CLKINVX1 U23 ( .A(n106), .Y(n11) );
  NAND2X1 U24 ( .A(n20), .B(n12), .Y(n122) );
  CLKINVX1 U25 ( .A(n86), .Y(n12) );
  CLKINVX1 U26 ( .A(n120), .Y(n4) );
  CLKINVX1 U27 ( .A(n119), .Y(n17) );
  CLKINVX1 U28 ( .A(n114), .Y(n5) );
  CLKINVX1 U29 ( .A(n107), .Y(n76) );
  NOR2X1 U30 ( .A(n20), .B(n7), .Y(n103) );
  NOR2X1 U31 ( .A(n16), .B(n7), .Y(n109) );
  INVX1 U32 ( .A(n125), .Y(n18) );
  AOI21X1 U33 ( .A0(n15), .A1(n7), .B0(n94), .Y(n120) );
  OAI21XL U34 ( .A0(n110), .A1(n130), .B0(n124), .Y(n82) );
  CLKINVX1 U36 ( .A(n81), .Y(n20) );
  NOR2X1 U37 ( .A(n18), .B(n13), .Y(n86) );
  NOR2X1 U38 ( .A(n124), .B(n107), .Y(n119) );
  OAI21XL U39 ( .A0(n109), .A1(n91), .B0(n130), .Y(n100) );
  NAND2X1 U40 ( .A(n103), .B(n87), .Y(n114) );
  CLKINVX1 U41 ( .A(n87), .Y(n14) );
  CLKINVX1 U42 ( .A(n91), .Y(n8) );
  CLKINVX1 U43 ( .A(n110), .Y(n9) );
  CLKINVX1 U44 ( .A(n121), .Y(n10) );
  OR2X1 U45 ( .A(n103), .B(n95), .Y(n126) );
  OAI221X1 U46 ( .A0(n18), .A1(n9), .B0(n7), .B1(n12), .C0(n93), .Y(n98) );
  AOI221XL U47 ( .A0(n95), .A1(n2), .B0(n92), .B1(n13), .C0(n6), .Y(n93) );
  OAI21XL U48 ( .A0(n1), .A1(n76), .B0(n8), .Y(n92) );
  XNOR2X1 U49 ( .A(addr[5]), .B(addr[3]), .Y(n102) );
  CLKINVX1 U51 ( .A(addr[5]), .Y(n77) );
  OAI221X1 U53 ( .A0(n76), .A1(n9), .B0(n16), .B1(n14), .C0(n105), .Y(n116) );
  AOI221XL U54 ( .A0(addr[3]), .A1(n104), .B0(n103), .B1(n130), .C0(n6), .Y(
        n105) );
  CLKINVX1 U55 ( .A(addr[6]), .Y(n78) );
  NAND3X1 U57 ( .A(n3), .B(n19), .C(n108), .Y(n113) );
  NOR2X1 U58 ( .A(n78), .B(addr[1]), .Y(n81) );
  AOI32XL U59 ( .A0(n1), .A1(n15), .A2(n124), .B0(n123), .B1(n78), .Y(n128) );
  AOI22XL U60 ( .A0(n2), .A1(n126), .B0(n125), .B1(n130), .Y(n127) );
  AOI222XL U61 ( .A0(n110), .A1(n125), .B0(n109), .B1(n15), .C0(n108), .C1(
        n107), .Y(n111) );
  OAI211XL U62 ( .A0(n106), .A1(n130), .B0(n1), .C0(addr[6]), .Y(n112) );
  OAI21XL U63 ( .A0(n3), .A1(addr[1]), .B0(n18), .Y(n80) );
  AOI221XL U64 ( .A0(n86), .A1(n15), .B0(n87), .B1(n125), .C0(n85), .Y(n89) );
  OAI211X1 U65 ( .A0(n84), .A1(n7), .B0(n83), .C0(n82), .Y(n85) );
  AOI222XL U66 ( .A0(n81), .A1(n15), .B0(n107), .B1(n106), .C0(n130), .C1(n19), 
        .Y(n84) );
  OAI21XL U67 ( .A0(n91), .A1(n6), .B0(addr[4]), .Y(n83) );
  AOI221XL U68 ( .A0(n125), .A1(n4), .B0(addr[3]), .B1(n126), .C0(n96), .Y(n97) );
  OAI22X1 U69 ( .A0(n16), .A1(n10), .B0(n11), .B1(n20), .Y(n96) );
  OAI211X1 U70 ( .A0(n76), .A1(n10), .B0(n118), .C0(n117), .Y(dout[3]) );
  AOI32XL U71 ( .A0(n125), .A1(n3), .A2(n102), .B0(n108), .B1(n109), .Y(n118)
         );
  AOI22XL U72 ( .A0(n116), .A1(n77), .B0(addr[5]), .B1(n115), .Y(n117) );
  AOI221XL U73 ( .A0(n121), .A1(n125), .B0(n95), .B1(n108), .C0(n5), .Y(n88)
         );
  AOI221XL U74 ( .A0(n130), .A1(n80), .B0(n94), .B1(n122), .C0(n79), .Y(n90)
         );
  NAND4X1 U75 ( .A(n101), .B(n113), .C(n100), .D(n99), .Y(dout[2]) );
  NAND3XL U76 ( .A(n2), .B(n124), .C(n102), .Y(n101) );
  AOI2BB2XL U77 ( .B0(addr[5]), .B1(n98), .A0N(addr[5]), .A1N(n97), .Y(n99) );
  OAI221X1 U78 ( .A0(n133), .A1(n77), .B0(n2), .B1(n132), .C0(n131), .Y(
        dout[4]) );
  AOI32XL U79 ( .A0(n130), .A1(n78), .A2(addr[2]), .B0(n129), .B1(n77), .Y(
        n131) );
  AOI222XL U80 ( .A0(n4), .A1(n122), .B0(n121), .B1(addr[1]), .C0(n120), .C1(
        n17), .Y(n133) );
  CLKINVX3 U81 ( .A(n2), .Y(n13) );
  CLKINVX3 U82 ( .A(addr[3]), .Y(n15) );
endmodule


module sbox4_7 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126;

  OAI32X4 U12 ( .A0(n16), .A1(n2), .A2(addr[2]), .B0(n72), .B1(n108), .Y(n123)
         );
  OAI222X4 U20 ( .A0(addr[2]), .A1(n92), .B0(n106), .B1(n91), .C0(n90), .C1(n9), .Y(dout[2]) );
  OAI222X4 U33 ( .A0(addr[4]), .A1(n106), .B0(n15), .B1(n108), .C0(n2), .C1(
        n118), .Y(n83) );
  NAND2X2 U34 ( .A(addr[4]), .B(n2), .Y(n108) );
  NOR2X2 U43 ( .A(n6), .B(addr[4]), .Y(n113) );
  NOR2X2 U45 ( .A(n72), .B(n2), .Y(n111) );
  NAND2X2 U51 ( .A(n15), .B(n12), .Y(n118) );
  NOR2X2 U52 ( .A(n71), .B(addr[5]), .Y(n97) );
  NAND2X2 U53 ( .A(addr[6]), .B(addr[1]), .Y(n85) );
  NAND2X2 U54 ( .A(addr[1]), .B(n12), .Y(n116) );
  NOR2X2 U55 ( .A(n115), .B(n72), .Y(n121) );
  NAND2X2 U56 ( .A(n6), .B(n71), .Y(n115) );
  NAND2X2 U57 ( .A(addr[5]), .B(n71), .Y(n96) );
  NAND2X2 U58 ( .A(addr[6]), .B(n15), .Y(n106) );
  OAI222X1 U1 ( .A0(n16), .A1(n85), .B0(n97), .B1(n116), .C0(n71), .C1(n118), 
        .Y(n73) );
  CLKINVX1 U2 ( .A(n116), .Y(n11) );
  CLKINVX1 U3 ( .A(n6), .Y(n1) );
  CLKBUFX3 U4 ( .A(addr[3]), .Y(n2) );
  OAI31X4 U5 ( .A0(n118), .A1(n72), .A2(n71), .B0(n117), .Y(n119) );
  OAI221X1 U6 ( .A0(addr[2]), .A1(n80), .B0(n118), .B1(n105), .C0(n79), .Y(
        dout[1]) );
  INVX4 U7 ( .A(addr[5]), .Y(n72) );
  OAI31X1 U8 ( .A0(n108), .A1(addr[5]), .A2(n13), .B0(n107), .Y(n109) );
  AOI222XL U9 ( .A0(n71), .A1(n12), .B0(n113), .B1(n15), .C0(addr[1]), .C1(n6), 
        .Y(n114) );
  OAI222X1 U10 ( .A0(addr[1]), .A1(n84), .B0(n85), .B1(n74), .C0(n6), .C1(n107), .Y(n75) );
  NAND2XL U11 ( .A(n1), .B(addr[5]), .Y(n84) );
  AOI211XL U13 ( .A0(n83), .A1(n72), .B0(n82), .C0(n5), .Y(n92) );
  NAND2XL U14 ( .A(n71), .B(n72), .Y(n74) );
  CLKINVX1 U15 ( .A(n118), .Y(n10) );
  CLKINVX1 U16 ( .A(n115), .Y(n4) );
  CLKINVX1 U17 ( .A(n112), .Y(n8) );
  OAI21X1 U18 ( .A0(n11), .A1(n13), .B0(n9), .Y(n112) );
  AOI22X1 U19 ( .A0(n14), .A1(n111), .B0(n13), .B1(n113), .Y(n93) );
  OAI211X1 U21 ( .A0(n15), .A1(n115), .B0(n93), .C0(n3), .Y(n94) );
  CLKINVX1 U22 ( .A(n85), .Y(n14) );
  NAND2X1 U23 ( .A(n97), .B(n6), .Y(n105) );
  NAND2X1 U24 ( .A(n113), .B(n10), .Y(n98) );
  NAND2X1 U25 ( .A(n11), .B(n97), .Y(n107) );
  NAND2X1 U26 ( .A(n118), .B(n85), .Y(n110) );
  OAI21XL U27 ( .A0(n4), .A1(n72), .B0(n108), .Y(n95) );
  CLKINVX1 U28 ( .A(n84), .Y(n7) );
  CLKINVX1 U29 ( .A(addr[2]), .Y(n9) );
  OAI31X1 U30 ( .A0(n71), .A1(addr[6]), .A2(n72), .B0(n87), .Y(n88) );
  OAI21XL U31 ( .A0(n113), .A1(n16), .B0(n14), .Y(n87) );
  OAI211X1 U32 ( .A0(n76), .A1(n71), .B0(n98), .C0(n3), .Y(n77) );
  AOI222XL U35 ( .A0(addr[5]), .A1(addr[6]), .B0(n111), .B1(addr[1]), .C0(n13), 
        .C1(n2), .Y(n76) );
  NAND3XL U36 ( .A(n14), .B(n6), .C(addr[4]), .Y(n117) );
  OAI22XL U37 ( .A0(n116), .A1(n115), .B0(n1), .B1(n112), .Y(n78) );
  CLKINVX3 U38 ( .A(addr[4]), .Y(n71) );
  OAI2BB2XL U39 ( .B0(n115), .B1(n106), .A0N(n72), .A1N(n86), .Y(n89) );
  OAI221XL U40 ( .A0(n116), .A1(addr[4]), .B0(n108), .B1(addr[1]), .C0(n117), 
        .Y(n86) );
  CLKINVX1 U41 ( .A(addr[6]), .Y(n12) );
  CLKINVX1 U42 ( .A(n81), .Y(n5) );
  OAI21XL U44 ( .A0(n96), .A1(n118), .B0(n93), .Y(n82) );
  NAND3X1 U46 ( .A(n101), .B(n100), .C(n99), .Y(n102) );
  AOI32X1 U47 ( .A0(n96), .A1(n6), .A2(n11), .B0(n14), .B1(n95), .Y(n101) );
  AOI2BB2XL U48 ( .B0(n15), .B1(n121), .A0N(n98), .A1N(addr[5]), .Y(n99) );
  OAI21XL U49 ( .A0(n97), .A1(n16), .B0(n13), .Y(n100) );
  AOI2BB2XL U50 ( .B0(n13), .B1(n123), .A0N(n122), .A1N(n9), .Y(n124) );
  AOI211XL U59 ( .A0(n13), .A1(n121), .B0(n120), .C0(n119), .Y(n122) );
  OAI22XL U60 ( .A0(n116), .A1(n115), .B0(addr[5]), .B1(n114), .Y(n120) );
  CLKINVX1 U61 ( .A(n75), .Y(n3) );
  AOI32XL U62 ( .A0(n11), .A1(n96), .A2(n1), .B0(addr[1]), .B1(n121), .Y(n81)
         );
  AOI222XL U63 ( .A0(n13), .A1(n16), .B0(n121), .B1(n116), .C0(n2), .C1(n73), 
        .Y(n80) );
  AOI22XL U64 ( .A0(n78), .A1(n72), .B0(addr[2]), .B1(n77), .Y(n79) );
  NAND2XL U65 ( .A(n111), .B(addr[4]), .Y(n91) );
  AOI211X1 U66 ( .A0(n7), .A1(n110), .B0(n89), .C0(n88), .Y(n90) );
  OAI211X1 U67 ( .A0(n106), .A1(n105), .B0(n104), .C0(n103), .Y(dout[3]) );
  AOI32X1 U68 ( .A0(n2), .A1(n16), .A2(n11), .B0(n94), .B1(n9), .Y(n104) );
  AOI22XL U69 ( .A0(addr[2]), .A1(n102), .B0(n10), .B1(n123), .Y(n103) );
  OAI211X1 U70 ( .A0(addr[2]), .A1(n126), .B0(n125), .C0(n124), .Y(dout[4]) );
  AOI32X1 U71 ( .A0(n14), .A1(n16), .A2(n2), .B0(n8), .B1(n7), .Y(n125) );
  AOI221XL U72 ( .A0(n10), .A1(n111), .B0(n4), .B1(n110), .C0(n109), .Y(n126)
         );
  CLKINVX3 U73 ( .A(n2), .Y(n6) );
  CLKINVX3 U74 ( .A(n106), .Y(n13) );
  CLKINVX3 U75 ( .A(addr[1]), .Y(n15) );
  CLKINVX3 U76 ( .A(n96), .Y(n16) );
endmodule


module sbox5_7 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121;

  OAI222X4 U18 ( .A0(addr[3]), .A1(n106), .B0(n8), .B1(n90), .C0(n13), .C1(n70), .Y(n93) );
  OAI22X2 U40 ( .A0(addr[5]), .A1(n106), .B0(n16), .B1(n114), .Y(n116) );
  NOR2X2 U41 ( .A(n3), .B(addr[3]), .Y(n102) );
  NAND2X2 U45 ( .A(addr[6]), .B(n70), .Y(n114) );
  NAND2X2 U50 ( .A(n70), .B(n8), .Y(n110) );
  NAND2X2 U52 ( .A(addr[1]), .B(n8), .Y(n113) );
  NAND2X2 U54 ( .A(addr[1]), .B(addr[6]), .Y(n106) );
  NAND2X2 U55 ( .A(addr[3]), .B(n13), .Y(n121) );
  CLKINVX1 U1 ( .A(addr[5]), .Y(n1) );
  AOI221XL U2 ( .A0(n93), .A1(n1), .B0(n9), .B1(n14), .C0(n92), .Y(n105) );
  INVX3 U3 ( .A(addr[5]), .Y(n16) );
  OAI221X4 U4 ( .A0(n111), .A1(n110), .B0(n121), .B1(n114), .C0(n109), .Y(n112) );
  OAI221X4 U5 ( .A0(n13), .A1(n114), .B0(n16), .B1(n113), .C0(n120), .Y(n115)
         );
  OAI221X4 U6 ( .A0(n107), .A1(n121), .B0(n111), .B1(n113), .C0(n85), .Y(n86)
         );
  OAI31X1 U7 ( .A0(n68), .A1(addr[5]), .A2(addr[1]), .B0(n81), .Y(n73) );
  OAI32X1 U8 ( .A0(n114), .A1(addr[5]), .A2(n3), .B0(n12), .B1(n107), .Y(n79)
         );
  AOI32XL U9 ( .A0(n14), .A1(n98), .A2(n7), .B0(n2), .B1(n73), .Y(n77) );
  CLKBUFX3 U10 ( .A(addr[4]), .Y(n2) );
  CLKINVX1 U11 ( .A(n81), .Y(n10) );
  NAND2X1 U12 ( .A(n11), .B(n14), .Y(n81) );
  CLKINVX1 U13 ( .A(n110), .Y(n5) );
  CLKXOR2X2 U14 ( .A(n68), .B(n16), .Y(n94) );
  AOI2BB1X1 U15 ( .A0N(n13), .A1N(n1), .B0(n14), .Y(n111) );
  NOR2X1 U16 ( .A(n121), .B(n16), .Y(n91) );
  NOR2BX1 U17 ( .AN(n116), .B(n90), .Y(n83) );
  NAND2X1 U19 ( .A(n5), .B(n16), .Y(n120) );
  CLKINVX1 U20 ( .A(n113), .Y(n7) );
  NAND2X1 U21 ( .A(n7), .B(n16), .Y(n107) );
  CLKINVX1 U22 ( .A(n121), .Y(n12) );
  OAI31X1 U23 ( .A0(n69), .A1(n14), .A2(n113), .B0(n99), .Y(n72) );
  CLKINVX1 U24 ( .A(n106), .Y(n9) );
  OAI2BB2XL U25 ( .B0(n1), .B1(n113), .A0N(n98), .A1N(n11), .Y(n101) );
  CLKINVX1 U26 ( .A(n114), .Y(n11) );
  CLKINVX1 U27 ( .A(n90), .Y(n15) );
  CLKINVX1 U28 ( .A(addr[1]), .Y(n70) );
  CLKINVX1 U29 ( .A(addr[3]), .Y(n68) );
  CLKINVX1 U30 ( .A(addr[6]), .Y(n8) );
  AOI211X1 U31 ( .A0(n91), .A1(addr[1]), .B0(n80), .C0(n79), .Y(n89) );
  OAI2BB2XL U32 ( .B0(n111), .B1(n106), .A0N(n94), .A1N(n5), .Y(n80) );
  AOI211X1 U33 ( .A0(n102), .A1(n84), .B0(n83), .C0(n82), .Y(n85) );
  OAI21XL U34 ( .A0(n8), .A1(n1), .B0(n106), .Y(n84) );
  NOR3XL U35 ( .A(n94), .B(n3), .C(n110), .Y(n82) );
  AOI222XL U36 ( .A0(n9), .A1(n15), .B0(addr[5]), .B1(n108), .C0(n6), .C1(n13), 
        .Y(n109) );
  CLKINVX1 U37 ( .A(n107), .Y(n6) );
  OAI21XL U38 ( .A0(addr[6]), .A1(addr[3]), .B0(n106), .Y(n108) );
  NAND2X1 U39 ( .A(addr[3]), .B(n3), .Y(n90) );
  NAND2X1 U42 ( .A(n2), .B(addr[5]), .Y(n98) );
  NAND2X1 U43 ( .A(n3), .B(n68), .Y(n97) );
  OAI21XL U44 ( .A0(addr[1]), .A1(n97), .B0(n96), .Y(n103) );
  AOI33XL U46 ( .A0(n3), .A1(n95), .A2(addr[5]), .B0(n94), .B1(n13), .B2(
        addr[1]), .Y(n96) );
  OAI21XL U47 ( .A0(n70), .A1(n68), .B0(n114), .Y(n95) );
  OAI21XL U48 ( .A0(addr[6]), .A1(n121), .B0(n99), .Y(n100) );
  NAND2X1 U49 ( .A(n71), .B(n5), .Y(n99) );
  XOR2X1 U51 ( .A(n69), .B(n3), .Y(n71) );
  AOI2BB2XL U53 ( .B0(n102), .B1(n116), .A0N(n2), .A1N(n75), .Y(n76) );
  AOI211X1 U56 ( .A0(n4), .A1(n3), .B0(n74), .C0(n83), .Y(n75) );
  AO22XL U57 ( .A0(n7), .A1(n12), .B0(addr[6]), .B1(n102), .Y(n74) );
  CLKINVX1 U58 ( .A(n120), .Y(n4) );
  CLKINVX1 U59 ( .A(n2), .Y(n69) );
  AO22XL U60 ( .A0(n7), .A1(n15), .B0(addr[6]), .B1(n91), .Y(n92) );
  AOI222XL U61 ( .A0(n116), .A1(n13), .B0(addr[3]), .B1(n115), .C0(n7), .C1(
        n14), .Y(n117) );
  OAI221X1 U62 ( .A0(n2), .A1(n105), .B0(n110), .B1(n121), .C0(n104), .Y(
        dout[3]) );
  AOI222XL U63 ( .A0(n2), .A1(n103), .B0(n102), .B1(n101), .C0(n100), .C1(n1), 
        .Y(n104) );
  OAI211X1 U64 ( .A0(n2), .A1(n89), .B0(n88), .C0(n87), .Y(dout[2]) );
  AOI33XL U65 ( .A0(n12), .A1(n98), .A2(n11), .B0(n3), .B1(n94), .B2(n5), .Y(
        n88) );
  AOI222XL U66 ( .A0(n10), .A1(n16), .B0(n2), .B1(n86), .C0(n91), .C1(n9), .Y(
        n87) );
  OAI211X1 U67 ( .A0(n78), .A1(n16), .B0(n77), .C0(n76), .Y(dout[1]) );
  AOI221XL U68 ( .A0(n12), .A1(addr[1]), .B0(n9), .B1(n14), .C0(n72), .Y(n78)
         );
  OAI211X1 U69 ( .A0(n121), .A1(n120), .B0(n119), .C0(n118), .Y(dout[4]) );
  AOI32XL U70 ( .A0(n14), .A1(n114), .A2(addr[5]), .B0(n2), .B1(n112), .Y(n119) );
  AOI2BB2X1 U71 ( .B0(n10), .B1(n16), .A0N(n2), .A1N(n117), .Y(n118) );
  BUFX4 U72 ( .A(addr[2]), .Y(n3) );
  CLKINVX3 U73 ( .A(n3), .Y(n13) );
  CLKINVX3 U74 ( .A(n97), .Y(n14) );
endmodule


module sbox6_7 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147;

  NAND2X2 U39 ( .A(n138), .B(addr[3]), .Y(n147) );
  NOR2X2 U47 ( .A(n7), .B(n17), .Y(n138) );
  NOR2X2 U50 ( .A(n13), .B(n4), .Y(n119) );
  NOR2X2 U58 ( .A(n84), .B(n13), .Y(n125) );
  NAND2X2 U61 ( .A(n97), .B(n103), .Y(n112) );
  NOR2X2 U62 ( .A(n85), .B(addr[1]), .Y(n103) );
  NOR2X2 U63 ( .A(n84), .B(addr[3]), .Y(n97) );
  NAND2X2 U64 ( .A(n117), .B(n131), .Y(n140) );
  NOR2X2 U65 ( .A(n5), .B(addr[3]), .Y(n131) );
  NOR2X2 U66 ( .A(n18), .B(addr[6]), .Y(n117) );
  NOR2X1 U1 ( .A(n7), .B(addr[3]), .Y(n102) );
  AOI211X1 U2 ( .A0(n15), .A1(n13), .B0(n131), .C0(n143), .Y(n121) );
  CLKINVX1 U3 ( .A(n84), .Y(n1) );
  INVX4 U4 ( .A(n4), .Y(n84) );
  CLKBUFX3 U5 ( .A(addr[4]), .Y(n4) );
  CLKINVX1 U6 ( .A(n7), .Y(n2) );
  OAI222X1 U7 ( .A0(n91), .A1(n15), .B0(n5), .B1(n14), .C0(addr[5]), .C1(n11), 
        .Y(n92) );
  BUFX4 U8 ( .A(addr[2]), .Y(n5) );
  OAI221X1 U9 ( .A0(n85), .A1(n12), .B0(n13), .B1(n16), .C0(n86), .Y(n90) );
  CLKINVX1 U10 ( .A(addr[3]), .Y(n3) );
  INVX3 U11 ( .A(addr[3]), .Y(n13) );
  OAI221X4 U12 ( .A0(n123), .A1(n82), .B0(n17), .B1(n15), .C0(n9), .Y(n124) );
  NOR2X4 U13 ( .A(addr[1]), .B(addr[6]), .Y(n130) );
  NOR2X4 U14 ( .A(n5), .B(addr[5]), .Y(n143) );
  INVX1 U15 ( .A(n130), .Y(n83) );
  CLKINVX1 U16 ( .A(n125), .Y(n12) );
  NAND2X1 U17 ( .A(n83), .B(n16), .Y(n105) );
  INVXL U18 ( .A(n121), .Y(n8) );
  CLKINVX1 U19 ( .A(n138), .Y(n6) );
  CLKINVX1 U20 ( .A(n117), .Y(n17) );
  CLKINVX1 U21 ( .A(n119), .Y(n11) );
  NOR2X1 U22 ( .A(n16), .B(n123), .Y(n144) );
  NOR2X1 U23 ( .A(n18), .B(n85), .Y(n96) );
  CLKINVX1 U24 ( .A(n103), .Y(n82) );
  OAI211X1 U25 ( .A0(n83), .A1(n12), .B0(n104), .C0(n112), .Y(n108) );
  OAI21XL U26 ( .A0(n103), .A1(n117), .B0(n102), .Y(n104) );
  OAI21XL U27 ( .A0(n132), .A1(n85), .B0(n3), .Y(n86) );
  AOI21X1 U28 ( .A0(n84), .A1(n102), .B0(n125), .Y(n91) );
  OAI2BB2XL U29 ( .B0(n143), .B1(n83), .A0N(n143), .A1N(n117), .Y(n118) );
  CLKINVX1 U30 ( .A(n122), .Y(n9) );
  CLKINVX1 U31 ( .A(n126), .Y(n81) );
  CLKINVX1 U32 ( .A(n97), .Y(n14) );
  NAND2BX1 U33 ( .AN(n144), .B(n137), .Y(n107) );
  CLKINVX1 U34 ( .A(addr[1]), .Y(n18) );
  NOR2X1 U35 ( .A(n16), .B(n2), .Y(n122) );
  NOR2X1 U36 ( .A(addr[1]), .B(n1), .Y(n132) );
  OAI22X1 U37 ( .A0(n11), .A1(n17), .B0(n5), .B1(n81), .Y(n88) );
  NAND2X1 U38 ( .A(n2), .B(n15), .Y(n123) );
  NAND4X1 U40 ( .A(n147), .B(n140), .C(n100), .D(n99), .Y(n101) );
  AOI222XL U41 ( .A0(n98), .A1(n7), .B0(n102), .B1(n130), .C0(n97), .C1(n105), 
        .Y(n99) );
  NAND3X1 U42 ( .A(n5), .B(n11), .C(n96), .Y(n100) );
  OAI221X1 U43 ( .A0(n13), .A1(n82), .B0(n11), .B1(n85), .C0(n81), .Y(n98) );
  AOI22X1 U44 ( .A0(n4), .A1(n115), .B0(addr[5]), .B1(n114), .Y(n129) );
  OAI21XL U45 ( .A0(n121), .A1(n83), .B0(n147), .Y(n115) );
  OAI21XL U46 ( .A0(n113), .A1(n7), .B0(n112), .Y(n114) );
  AOI221XL U48 ( .A0(n119), .A1(n18), .B0(n130), .B1(addr[3]), .C0(n111), .Y(
        n113) );
  OAI22XL U49 ( .A0(n17), .A1(n84), .B0(addr[3]), .B1(n16), .Y(n111) );
  OAI22XL U51 ( .A0(n13), .A1(n85), .B0(addr[1]), .B1(n11), .Y(n142) );
  AOI211X1 U52 ( .A0(n4), .A1(n135), .B0(n134), .C0(n133), .Y(n136) );
  OA21XL U53 ( .A0(n3), .A1(n2), .B0(n132), .Y(n133) );
  OAI2BB2XL U54 ( .B0(n1), .B1(n9), .A0N(n131), .A1N(n130), .Y(n134) );
  OAI22X1 U55 ( .A0(n5), .A1(n17), .B0(n7), .B1(n16), .Y(n135) );
  CLKINVX3 U56 ( .A(addr[5]), .Y(n15) );
  AOI2BB2X1 U57 ( .B0(n5), .B1(n130), .A0N(n2), .A1N(n82), .Y(n137) );
  NOR2X1 U59 ( .A(n82), .B(n1), .Y(n126) );
  AOI2BB2XL U60 ( .B0(n143), .B1(n90), .A0N(n89), .A1N(n15), .Y(n94) );
  AOI211X1 U67 ( .A0(n122), .A1(n4), .B0(n88), .C0(n87), .Y(n89) );
  OAI32X1 U68 ( .A0(n82), .A1(n13), .A2(n7), .B0(n6), .B1(n14), .Y(n87) );
  NAND3X1 U69 ( .A(n147), .B(n140), .C(n139), .Y(n141) );
  AOI32X1 U70 ( .A0(n5), .A1(n18), .A2(n4), .B0(n138), .B1(n84), .Y(n139) );
  AO22XL U71 ( .A0(n143), .A1(n1), .B0(n116), .B1(n84), .Y(n120) );
  OAI21XL U72 ( .A0(n2), .A1(n15), .B0(n123), .Y(n116) );
  CLKINVX1 U73 ( .A(n106), .Y(n10) );
  AOI32XL U74 ( .A0(n105), .A1(n84), .A2(n3), .B0(addr[1]), .B1(n125), .Y(n106) );
  OAI211X1 U75 ( .A0(n84), .A1(n140), .B0(n110), .C0(n109), .Y(dout[2]) );
  AOI222XL U76 ( .A0(n108), .A1(n15), .B0(n143), .B1(n10), .C0(n119), .C1(n107), .Y(n109) );
  AOI2BB2XL U77 ( .B0(addr[5]), .B1(n101), .A0N(n7), .A1N(n112), .Y(n110) );
  OAI211X1 U78 ( .A0(n1), .A1(n147), .B0(n146), .C0(n145), .Y(dout[4]) );
  AOI222XL U79 ( .A0(n144), .A1(n13), .B0(n143), .B1(n142), .C0(n141), .C1(n15), .Y(n145) );
  OA22X1 U80 ( .A0(n12), .A1(n137), .B0(n136), .B1(n15), .Y(n146) );
  NAND3X1 U81 ( .A(n129), .B(n128), .C(n127), .Y(dout[3]) );
  AOI32XL U82 ( .A0(n120), .A1(n13), .A2(addr[1]), .B0(n119), .B1(n118), .Y(
        n128) );
  AOI222XL U83 ( .A0(n144), .A1(n84), .B0(n126), .B1(n8), .C0(n125), .C1(n124), 
        .Y(n127) );
  NAND3BX1 U84 ( .AN(n95), .B(n94), .C(n93), .Y(dout[1]) );
  OAI222X1 U85 ( .A0(n140), .A1(n4), .B0(n112), .B1(n7), .C0(n16), .C1(n91), 
        .Y(n95) );
  AOI32XL U86 ( .A0(addr[1]), .A1(n15), .A2(n125), .B0(n130), .B1(n92), .Y(n93) );
  CLKINVX3 U87 ( .A(n5), .Y(n7) );
  CLKINVX3 U88 ( .A(n96), .Y(n16) );
  CLKINVX3 U89 ( .A(addr[6]), .Y(n85) );
endmodule


module sbox7_7 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148;

  OAI222X4 U19 ( .A0(n11), .A1(n129), .B0(n4), .B1(n7), .C0(addr[1]), .C1(n18), 
        .Y(n122) );
  OAI33X4 U33 ( .A0(addr[1]), .A1(n4), .A2(n5), .B0(n8), .B1(n86), .B2(n12), 
        .Y(n97) );
  NOR2X2 U44 ( .A(n16), .B(n4), .Y(n116) );
  NOR2X2 U48 ( .A(addr[1]), .B(addr[6]), .Y(n136) );
  NOR2X2 U51 ( .A(n21), .B(n16), .Y(n125) );
  NOR2X2 U52 ( .A(n8), .B(addr[3]), .Y(n131) );
  NOR2X2 U58 ( .A(n93), .B(n124), .Y(n142) );
  NOR2X2 U60 ( .A(n85), .B(addr[1]), .Y(n93) );
  NOR2X2 U62 ( .A(n87), .B(n3), .Y(n137) );
  NOR2X2 U65 ( .A(n85), .B(n9), .Y(n140) );
  NAND2X1 U1 ( .A(n3), .B(n4), .Y(n119) );
  CLKBUFX3 U2 ( .A(addr[4]), .Y(n4) );
  CLKINVX1 U3 ( .A(n87), .Y(n1) );
  CLKINVX1 U4 ( .A(n86), .Y(n2) );
  CLKBUFX3 U5 ( .A(addr[2]), .Y(n5) );
  OAI22X1 U6 ( .A0(addr[1]), .A1(n18), .B0(n5), .B1(n113), .Y(n100) );
  OAI31X1 U7 ( .A0(n16), .A1(n87), .A2(n9), .B0(n117), .Y(n121) );
  OAI22X1 U8 ( .A0(n4), .A1(n21), .B0(addr[3]), .B1(n84), .Y(n103) );
  NOR2X4 U9 ( .A(n9), .B(addr[6]), .Y(n124) );
  AOI211XL U10 ( .A0(n5), .A1(n6), .B0(n131), .C0(n130), .Y(n132) );
  NOR3XL U11 ( .A(n11), .B(addr[3]), .C(n2), .Y(n130) );
  OAI21XL U12 ( .A0(n3), .A1(n1), .B0(n119), .Y(n89) );
  BUFX4 U13 ( .A(addr[5]), .Y(n3) );
  AOI221XL U14 ( .A0(n140), .A1(n89), .B0(n109), .B1(n6), .C0(n88), .Y(n96) );
  CLKINVX1 U15 ( .A(n140), .Y(n8) );
  OAI2BB2XL U16 ( .B0(n142), .B1(n84), .A0N(n141), .A1N(n140), .Y(n143) );
  CLKINVX1 U17 ( .A(n125), .Y(n14) );
  CLKINVX1 U18 ( .A(n142), .Y(n6) );
  NAND2X1 U20 ( .A(n14), .B(n19), .Y(n105) );
  CLKINVX1 U21 ( .A(n123), .Y(n17) );
  CLKINVX1 U22 ( .A(n109), .Y(n15) );
  NAND2X1 U23 ( .A(n124), .B(n16), .Y(n113) );
  CLKINVX1 U24 ( .A(n137), .Y(n84) );
  NOR2X1 U25 ( .A(n84), .B(n16), .Y(n109) );
  CLKINVX1 U26 ( .A(n136), .Y(n11) );
  OAI22XL U27 ( .A0(n137), .A1(n7), .B0(n9), .B1(n15), .Y(n146) );
  OAI21X1 U28 ( .A0(n87), .A1(n14), .B0(n129), .Y(n141) );
  NAND2X1 U29 ( .A(n116), .B(n21), .Y(n129) );
  CLKINVX1 U30 ( .A(n93), .Y(n10) );
  OAI21XL U31 ( .A0(n119), .A1(n10), .B0(n118), .Y(n120) );
  OAI21XL U32 ( .A0(n125), .A1(n137), .B0(n124), .Y(n118) );
  NOR2X1 U34 ( .A(n21), .B(n18), .Y(n123) );
  CLKINVX1 U35 ( .A(n145), .Y(n18) );
  OAI22XL U36 ( .A0(n137), .A1(n113), .B0(n85), .B1(n17), .Y(n88) );
  CLKINVX1 U37 ( .A(n116), .Y(n12) );
  CLKINVX1 U38 ( .A(n131), .Y(n7) );
  CLKINVX1 U39 ( .A(n134), .Y(n19) );
  NOR2XL U40 ( .A(n125), .B(n87), .Y(n110) );
  CLKINVX1 U41 ( .A(n119), .Y(n83) );
  CLKINVX1 U42 ( .A(n103), .Y(n20) );
  OA21XL U43 ( .A0(n13), .A1(n10), .B0(n117), .Y(n102) );
  CLKINVX1 U45 ( .A(n105), .Y(n13) );
  OAI2BB1XL U46 ( .A0N(n103), .A1N(n124), .B0(n102), .Y(n104) );
  OAI22X1 U47 ( .A0(n21), .A1(n12), .B0(n4), .B1(n19), .Y(n112) );
  NOR4X1 U49 ( .A(n4), .B(addr[3]), .C(n9), .D(n86), .Y(n99) );
  XNOR2X1 U50 ( .A(addr[6]), .B(n5), .Y(n101) );
  AOI211X1 U53 ( .A0(n116), .A1(addr[6]), .B0(n115), .C0(n114), .Y(n128) );
  OAI222X1 U54 ( .A0(n111), .A1(n8), .B0(n110), .B1(n10), .C0(n11), .C1(n15), 
        .Y(n115) );
  OAI2BB2XL U55 ( .B0(n83), .B1(n113), .A0N(n9), .A1N(n112), .Y(n114) );
  OA21XL U56 ( .A0(n16), .A1(n3), .B0(n17), .Y(n111) );
  NAND2X1 U57 ( .A(n5), .B(n136), .Y(n133) );
  CLKINVX1 U59 ( .A(addr[6]), .Y(n85) );
  AOI211X1 U61 ( .A0(n131), .A1(n3), .B0(n92), .C0(n91), .Y(n95) );
  OAI221X1 U63 ( .A0(n9), .A1(n18), .B0(n8), .B1(n84), .C0(n102), .Y(n92) );
  OAI31X1 U64 ( .A0(n16), .A1(n87), .A2(n11), .B0(n90), .Y(n91) );
  AO21XL U66 ( .A0(n119), .A1(n129), .B0(addr[6]), .Y(n90) );
  NOR2X1 U67 ( .A(n87), .B(addr[3]), .Y(n145) );
  AOI21XL U68 ( .A0(addr[3]), .A1(n98), .B0(n97), .Y(n108) );
  OAI2BB1XL U69 ( .A0N(n86), .A1N(n124), .B0(n133), .Y(n98) );
  NAND3X1 U70 ( .A(n136), .B(n16), .C(n3), .Y(n117) );
  NOR2X1 U71 ( .A(addr[3]), .B(n3), .Y(n134) );
  OAI21X1 U72 ( .A0(n5), .A1(n142), .B0(n133), .Y(n138) );
  OAI22XL U73 ( .A0(n142), .A1(n12), .B0(n1), .B1(n132), .Y(n135) );
  AO21X1 U74 ( .A0(n139), .A1(n21), .B0(n138), .Y(n144) );
  OAI21XL U75 ( .A0(n2), .A1(n9), .B0(n10), .Y(n139) );
  OAI221X1 U76 ( .A0(n96), .A1(n86), .B0(n5), .B1(n95), .C0(n94), .Y(dout[1])
         );
  AOI2BB2X1 U77 ( .B0(n93), .B1(n112), .A0N(n133), .A1N(n20), .Y(n94) );
  OAI211X1 U78 ( .A0(n128), .A1(n86), .B0(n127), .C0(n126), .Y(dout[3]) );
  AOI32XL U79 ( .A0(n125), .A1(n1), .A2(n124), .B0(n123), .B1(n136), .Y(n126)
         );
  OAI31X1 U80 ( .A0(n122), .A1(n121), .A2(n120), .B0(n86), .Y(n127) );
  OAI221X1 U81 ( .A0(n3), .A1(n108), .B0(n107), .B1(n21), .C0(n106), .Y(
        dout[2]) );
  AOI32XL U82 ( .A0(n105), .A1(n86), .A2(n140), .B0(n2), .B1(n104), .Y(n106)
         );
  AOI211X1 U83 ( .A0(n101), .A1(n4), .B0(n100), .C0(n99), .Y(n107) );
  NAND2X1 U84 ( .A(n148), .B(n147), .Y(dout[4]) );
  AOI222XL U85 ( .A0(n136), .A1(n141), .B0(n3), .B1(n135), .C0(n134), .C1(n138), .Y(n148) );
  AOI222XL U86 ( .A0(n5), .A1(n146), .B0(n145), .B1(n144), .C0(n143), .C1(n86), 
        .Y(n147) );
  CLKINVX3 U87 ( .A(addr[1]), .Y(n9) );
  CLKINVX3 U88 ( .A(addr[3]), .Y(n16) );
  CLKINVX3 U89 ( .A(n3), .Y(n21) );
  CLKINVX3 U90 ( .A(n5), .Y(n86) );
  CLKINVX3 U91 ( .A(n4), .Y(n87) );
endmodule


module sbox8_7 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132;

  NAND2X2 U41 ( .A(addr[6]), .B(n10), .Y(n131) );
  NAND2X2 U48 ( .A(addr[4]), .B(n16), .Y(n123) );
  NAND2X2 U49 ( .A(n2), .B(n74), .Y(n87) );
  NAND2X2 U50 ( .A(addr[1]), .B(n6), .Y(n124) );
  NAND2X2 U54 ( .A(addr[2]), .B(n75), .Y(n116) );
  NAND2X2 U60 ( .A(addr[6]), .B(addr[1]), .Y(n105) );
  NAND2X2 U61 ( .A(n10), .B(n6), .Y(n108) );
  OAI32X1 U1 ( .A0(n6), .A1(addr[4]), .A2(n92), .B0(n115), .B1(n108), .Y(n96)
         );
  OAI31X1 U2 ( .A0(n123), .A1(addr[6]), .A2(n116), .B0(n109), .Y(n110) );
  AOI222X1 U3 ( .A0(n88), .A1(addr[2]), .B0(n74), .B1(n11), .C0(n12), .C1(n92), 
        .Y(n114) );
  OAI222X1 U4 ( .A0(addr[2]), .A1(n126), .B0(n16), .B1(n125), .C0(n124), .C1(
        n123), .Y(n127) );
  OAI221X1 U5 ( .A0(n105), .A1(n87), .B0(addr[4]), .B1(n108), .C0(n86), .Y(n90) );
  NAND2X4 U6 ( .A(addr[4]), .B(n2), .Y(n115) );
  AOI32XL U7 ( .A0(n4), .A1(n14), .A2(n2), .B0(n5), .B1(n117), .Y(n130) );
  OA21XL U8 ( .A0(n12), .A1(n75), .B0(n121), .Y(n78) );
  INVXL U9 ( .A(n119), .Y(n3) );
  INVX3 U10 ( .A(n2), .Y(n16) );
  BUFX4 U11 ( .A(addr[3]), .Y(n2) );
  CLKBUFX3 U12 ( .A(addr[5]), .Y(n1) );
  CLKINVX1 U13 ( .A(n108), .Y(n5) );
  CLKINVX1 U14 ( .A(n107), .Y(n13) );
  CLKINVX1 U15 ( .A(n93), .Y(n15) );
  NAND2X1 U16 ( .A(n16), .B(n74), .Y(n93) );
  NAND2X1 U17 ( .A(n12), .B(n75), .Y(n121) );
  OAI21XL U18 ( .A0(n115), .A1(n75), .B0(n107), .Y(n77) );
  OAI21X1 U19 ( .A0(n74), .A1(n75), .B0(n123), .Y(n88) );
  OAI31XL U20 ( .A0(n115), .A1(n10), .A2(n116), .B0(n118), .Y(n94) );
  CLKINVX1 U21 ( .A(n131), .Y(n9) );
  NAND2X1 U22 ( .A(n14), .B(n16), .Y(n107) );
  OAI22XL U23 ( .A0(n116), .A1(n123), .B0(n14), .B1(n115), .Y(n117) );
  OAI22XL U24 ( .A0(n123), .A1(n108), .B0(n131), .B1(n93), .Y(n95) );
  OAI2BB2XL U25 ( .B0(n115), .B1(n131), .A0N(n88), .A1N(n8), .Y(n89) );
  AOI211XL U26 ( .A0(n108), .A1(n105), .B0(n74), .C0(n121), .Y(n85) );
  CLKINVX1 U27 ( .A(n124), .Y(n4) );
  OAI22XL U28 ( .A0(n14), .A1(n123), .B0(n78), .B1(n87), .Y(n81) );
  NAND2BX2 U29 ( .AN(n78), .B(n16), .Y(n120) );
  NAND2XL U30 ( .A(n115), .B(n93), .Y(n104) );
  OAI2BB2XL U31 ( .B0(n106), .B1(n105), .A0N(n104), .A1N(n4), .Y(n111) );
  NOR2BXL U32 ( .AN(n123), .B(n103), .Y(n106) );
  NAND3X1 U33 ( .A(n104), .B(n10), .C(n14), .Y(n84) );
  AO21X1 U34 ( .A0(n14), .A1(n8), .B0(n101), .Y(n102) );
  OAI33X1 U35 ( .A0(n6), .A1(n16), .A2(n100), .B0(n12), .B1(n103), .B2(n124), 
        .Y(n101) );
  OA22XL U36 ( .A0(n107), .A1(n131), .B0(n120), .B1(n124), .Y(n98) );
  CLKINVX1 U37 ( .A(n125), .Y(n7) );
  OAI21XL U38 ( .A0(n4), .A1(n9), .B0(addr[4]), .Y(n86) );
  NAND2X1 U39 ( .A(n1), .B(n12), .Y(n100) );
  OAI221X1 U40 ( .A0(n124), .A1(n121), .B0(addr[1]), .B1(n120), .C0(n3), .Y(
        n128) );
  OAI31XL U42 ( .A0(n12), .A1(n10), .A2(n16), .B0(n118), .Y(n119) );
  NAND2X1 U43 ( .A(n8), .B(addr[2]), .Y(n125) );
  NAND4XL U44 ( .A(n9), .B(n1), .C(n2), .D(addr[2]), .Y(n109) );
  NAND3X1 U45 ( .A(n14), .B(n6), .C(n2), .Y(n118) );
  OAI21XL U46 ( .A0(n1), .A1(n87), .B0(n114), .Y(n76) );
  OAI22XL U47 ( .A0(n108), .A1(n120), .B0(n79), .B1(n100), .Y(n80) );
  AOI221XL U51 ( .A0(n9), .A1(n16), .B0(n8), .B1(n2), .C0(n91), .Y(n79) );
  NOR2X1 U52 ( .A(n1), .B(n2), .Y(n103) );
  NOR2X1 U53 ( .A(n87), .B(addr[6]), .Y(n91) );
  NOR2X1 U55 ( .A(n16), .B(n1), .Y(n92) );
  CLKINVX1 U56 ( .A(n100), .Y(n11) );
  OA21XL U57 ( .A0(n1), .A1(n115), .B0(n120), .Y(n132) );
  AOI221XL U58 ( .A0(n5), .A1(n2), .B0(n8), .B1(addr[4]), .C0(n122), .Y(n126)
         );
  OAI22XL U59 ( .A0(n2), .A1(n10), .B0(addr[4]), .B1(n131), .Y(n122) );
  OAI211X1 U62 ( .A0(addr[2]), .A1(n99), .B0(n98), .C0(n97), .Y(dout[2]) );
  AOI221XL U63 ( .A0(addr[2]), .A1(n96), .B0(n1), .B1(n95), .C0(n94), .Y(n97)
         );
  AOI221XL U64 ( .A0(n91), .A1(n1), .B0(n90), .B1(n75), .C0(n89), .Y(n99) );
  OAI211X1 U65 ( .A0(n132), .A1(n131), .B0(n130), .C0(n129), .Y(dout[4]) );
  AOI222XL U66 ( .A0(n128), .A1(n74), .B0(n1), .B1(n127), .C0(n13), .C1(n8), 
        .Y(n129) );
  OAI211X1 U67 ( .A0(addr[1]), .A1(n114), .B0(n113), .C0(n112), .Y(dout[3]) );
  AOI221XL U68 ( .A0(n111), .A1(n12), .B0(n13), .B1(n5), .C0(n110), .Y(n112)
         );
  AOI2BB2XL U69 ( .B0(n102), .B1(n74), .A0N(n115), .A1N(n125), .Y(n113) );
  NAND4BX1 U70 ( .AN(n85), .B(n84), .C(n83), .D(n82), .Y(dout[1]) );
  AOI221XL U71 ( .A0(n9), .A1(n81), .B0(n15), .B1(n7), .C0(n80), .Y(n82) );
  AOI22X1 U72 ( .A0(n8), .A1(n77), .B0(n4), .B1(n76), .Y(n83) );
  CLKINVX3 U73 ( .A(addr[6]), .Y(n6) );
  CLKINVX3 U74 ( .A(n105), .Y(n8) );
  CLKINVX3 U75 ( .A(addr[1]), .Y(n10) );
  CLKINVX3 U76 ( .A(addr[2]), .Y(n12) );
  CLKINVX3 U77 ( .A(n116), .Y(n14) );
  CLKINVX3 U78 ( .A(addr[4]), .Y(n74) );
  CLKINVX3 U79 ( .A(n1), .Y(n75) );
endmodule


module crp_7 ( P, R, K_sub );
  output [1:32] P;
  input [1:32] R;
  input [1:48] K_sub;
  wire   n1;
  wire   [1:48] X;

  sbox1_7 u0 ( .addr(X[1:6]), .dout({P[9], P[17], P[23], P[31]}) );
  sbox2_7 u1 ( .addr({X[7], n1, X[9:12]}), .dout({P[13], P[28], P[2], P[18]})
         );
  sbox3_7 u2 ( .addr(X[13:18]), .dout({P[24], P[16], P[30], P[6]}) );
  sbox4_7 u3 ( .addr(X[19:24]), .dout({P[26], P[20], P[10], P[1]}) );
  sbox5_7 u4 ( .addr(X[25:30]), .dout({P[8], P[14], P[25], P[3]}) );
  sbox6_7 u5 ( .addr(X[31:36]), .dout({P[4], P[29], P[11], P[19]}) );
  sbox7_7 u6 ( .addr(X[37:42]), .dout({P[32], P[12], P[22], P[7]}) );
  sbox8_7 u7 ( .addr(X[43:48]), .dout({P[5], P[27], P[15], P[21]}) );
  XOR2X1 U1 ( .A(R[1]), .B(K_sub[2]), .Y(X[2]) );
  CLKXOR2X4 U2 ( .A(R[29]), .B(K_sub[42]), .Y(X[42]) );
  CLKXOR2X4 U3 ( .A(R[5]), .B(K_sub[6]), .Y(X[6]) );
  CLKXOR2X4 U4 ( .A(R[16]), .B(K_sub[25]), .Y(X[25]) );
  CLKXOR2X4 U5 ( .A(R[29]), .B(K_sub[44]), .Y(X[44]) );
  CLKXOR2X4 U6 ( .A(R[22]), .B(K_sub[33]), .Y(X[33]) );
  CLKXOR2X4 U7 ( .A(R[8]), .B(K_sub[11]), .Y(X[11]) );
  CLKXOR2X4 U8 ( .A(R[16]), .B(K_sub[23]), .Y(X[23]) );
  CLKXOR2X4 U9 ( .A(R[26]), .B(K_sub[39]), .Y(X[39]) );
  CLKXOR2X4 U10 ( .A(R[10]), .B(K_sub[15]), .Y(X[15]) );
  XNOR2X1 U11 ( .A(R[5]), .B(K_sub[8]), .Y(X[8]) );
  INVX3 U12 ( .A(X[8]), .Y(n1) );
  CLKXOR2X4 U13 ( .A(R[20]), .B(K_sub[31]), .Y(X[31]) );
  CLKXOR2X4 U14 ( .A(R[31]), .B(K_sub[46]), .Y(X[46]) );
  CLKXOR2X4 U15 ( .A(R[12]), .B(K_sub[19]), .Y(X[19]) );
  CLKXOR2X4 U16 ( .A(R[20]), .B(K_sub[29]), .Y(X[29]) );
  CLKXOR2X2 U17 ( .A(R[4]), .B(K_sub[5]), .Y(X[5]) );
  CLKXOR2X2 U18 ( .A(R[15]), .B(K_sub[22]), .Y(X[22]) );
  CLKXOR2X2 U19 ( .A(R[24]), .B(K_sub[35]), .Y(X[35]) );
  CLKXOR2X2 U20 ( .A(R[21]), .B(K_sub[30]), .Y(X[30]) );
  CLKXOR2X2 U21 ( .A(R[12]), .B(K_sub[17]), .Y(X[17]) );
  CLKXOR2X2 U22 ( .A(R[32]), .B(K_sub[1]), .Y(X[1]) );
  CLKXOR2X2 U23 ( .A(R[13]), .B(K_sub[20]), .Y(X[20]) );
  CLKXOR2X2 U24 ( .A(R[18]), .B(K_sub[27]), .Y(X[27]) );
  CLKXOR2X2 U25 ( .A(R[8]), .B(K_sub[13]), .Y(X[13]) );
  CLKXOR2X2 U26 ( .A(R[4]), .B(K_sub[7]), .Y(X[7]) );
  CLKXOR2X2 U27 ( .A(R[24]), .B(K_sub[37]), .Y(X[37]) );
  CLKXOR2X2 U28 ( .A(R[28]), .B(K_sub[43]), .Y(X[43]) );
  CLKXOR2X2 U29 ( .A(R[1]), .B(K_sub[48]), .Y(X[48]) );
  CLKXOR2X2 U30 ( .A(R[17]), .B(K_sub[24]), .Y(X[24]) );
  CLKXOR2X2 U31 ( .A(R[9]), .B(K_sub[12]), .Y(X[12]) );
  CLKXOR2X2 U32 ( .A(R[13]), .B(K_sub[18]), .Y(X[18]) );
  CLKXOR2X2 U33 ( .A(R[25]), .B(K_sub[36]), .Y(X[36]) );
  XOR2X1 U34 ( .A(R[23]), .B(K_sub[34]), .Y(X[34]) );
  XOR2X1 U35 ( .A(R[9]), .B(K_sub[14]), .Y(X[14]) );
  XOR2X1 U36 ( .A(R[30]), .B(K_sub[45]), .Y(X[45]) );
  XOR2X1 U37 ( .A(R[21]), .B(K_sub[32]), .Y(X[32]) );
  XOR2X1 U38 ( .A(R[25]), .B(K_sub[38]), .Y(X[38]) );
  XOR2X1 U39 ( .A(R[27]), .B(K_sub[40]), .Y(X[40]) );
  XOR2X1 U40 ( .A(R[3]), .B(K_sub[4]), .Y(X[4]) );
  XOR2X1 U41 ( .A(R[11]), .B(K_sub[16]), .Y(X[16]) );
  XOR2X1 U42 ( .A(R[7]), .B(K_sub[10]), .Y(X[10]) );
  XOR2X1 U43 ( .A(R[14]), .B(K_sub[21]), .Y(X[21]) );
  XOR2X1 U44 ( .A(R[6]), .B(K_sub[9]), .Y(X[9]) );
  XOR2X1 U45 ( .A(R[2]), .B(K_sub[3]), .Y(X[3]) );
  XOR2X1 U46 ( .A(R[28]), .B(K_sub[41]), .Y(X[41]) );
  XOR2X1 U47 ( .A(R[17]), .B(K_sub[26]), .Y(X[26]) );
  XOR2X1 U48 ( .A(R[32]), .B(K_sub[47]), .Y(X[47]) );
  XOR2X1 U49 ( .A(R[19]), .B(K_sub[28]), .Y(X[28]) );
endmodule


module sbox1_6 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127;

  OAI222X4 U13 ( .A0(addr[5]), .A1(n101), .B0(n1), .B1(n100), .C0(n99), .C1(n6), .Y(dout[3]) );
  OAI21X2 U42 ( .A0(n4), .A1(n112), .B0(n106), .Y(n123) );
  NAND2X2 U44 ( .A(addr[6]), .B(n10), .Y(n115) );
  NAND2X2 U48 ( .A(addr[1]), .B(n13), .Y(n114) );
  OAI22X2 U49 ( .A0(n69), .A1(n72), .B0(addr[5]), .B1(n120), .Y(n85) );
  NAND2X2 U50 ( .A(n3), .B(n69), .Y(n120) );
  NOR2X2 U51 ( .A(n69), .B(n3), .Y(n124) );
  NOR2X2 U56 ( .A(n109), .B(n3), .Y(n93) );
  NAND2X2 U57 ( .A(addr[1]), .B(addr[6]), .Y(n109) );
  NAND2X2 U59 ( .A(n10), .B(n13), .Y(n112) );
  NOR2X1 U1 ( .A(n114), .B(n120), .Y(n104) );
  AOI221X4 U2 ( .A0(n9), .A1(n90), .B0(n4), .B1(n93), .C0(n102), .Y(n79) );
  NOR3X1 U3 ( .A(n2), .B(addr[6]), .C(n6), .Y(n102) );
  BUFX4 U4 ( .A(addr[4]), .Y(n2) );
  CLKBUFX3 U5 ( .A(addr[2]), .Y(n1) );
  OAI32X1 U6 ( .A0(n112), .A1(n2), .A2(n4), .B0(n115), .B1(n113), .Y(n80) );
  NOR2BXL U7 ( .AN(n118), .B(n1), .Y(n122) );
  CLKBUFX3 U8 ( .A(addr[2]), .Y(n4) );
  OAI221X4 U9 ( .A0(addr[5]), .A1(n127), .B0(n126), .B1(n72), .C0(n125), .Y(
        dout[4]) );
  OAI221X4 U10 ( .A0(n88), .A1(n72), .B0(addr[5]), .B1(n87), .C0(n86), .Y(
        dout[2]) );
  OA21XL U11 ( .A0(n95), .A1(n115), .B0(n107), .Y(n119) );
  AOI222XL U12 ( .A0(n9), .A1(n1), .B0(n2), .B1(n110), .C0(n11), .C1(n6), .Y(
        n111) );
  AOI2BB2X1 U14 ( .B0(n2), .B1(n11), .A0N(addr[4]), .A1N(n115), .Y(n91) );
  BUFX4 U15 ( .A(addr[3]), .Y(n3) );
  CLKINVX1 U16 ( .A(n112), .Y(n9) );
  CLKINVX1 U17 ( .A(n113), .Y(n5) );
  NAND2BX1 U18 ( .AN(n104), .B(n119), .Y(n84) );
  CLKXOR2X2 U19 ( .A(n70), .B(n6), .Y(n90) );
  NOR2X1 U20 ( .A(n69), .B(n70), .Y(n118) );
  OAI21XL U21 ( .A0(n70), .A1(n114), .B0(n91), .Y(n92) );
  NAND2X1 U22 ( .A(n93), .B(n69), .Y(n107) );
  NAND2X1 U23 ( .A(n6), .B(n70), .Y(n113) );
  OAI211X1 U24 ( .A0(n69), .A1(n114), .B0(n108), .C0(n107), .Y(n89) );
  CLKINVX1 U25 ( .A(n109), .Y(n11) );
  NAND2X1 U26 ( .A(n124), .B(n8), .Y(n108) );
  CLKINVX1 U27 ( .A(n114), .Y(n12) );
  CLKINVX1 U28 ( .A(n115), .Y(n8) );
  CLKINVX1 U29 ( .A(n95), .Y(n71) );
  AO22X1 U30 ( .A0(n90), .A1(n8), .B0(n70), .B1(n123), .Y(n76) );
  OAI31X1 U31 ( .A0(n6), .A1(n3), .A2(n10), .B0(n103), .Y(n105) );
  AOI31XL U32 ( .A0(n10), .A1(n6), .A2(n2), .B0(n102), .Y(n103) );
  CLKINVX1 U33 ( .A(addr[6]), .Y(n13) );
  AOI211X1 U34 ( .A0(n7), .A1(n4), .B0(n117), .C0(n116), .Y(n126) );
  CLKINVX1 U35 ( .A(n108), .Y(n7) );
  AOI211X1 U36 ( .A0(n115), .A1(n114), .B0(n113), .C0(n2), .Y(n116) );
  OAI22X1 U37 ( .A0(n120), .A1(n112), .B0(n111), .B1(n70), .Y(n117) );
  AOI211X1 U38 ( .A0(n11), .A1(n118), .B0(n81), .C0(n80), .Y(n88) );
  OAI22X1 U39 ( .A0(n91), .A1(n6), .B0(n3), .B1(n106), .Y(n81) );
  CLKINVX3 U40 ( .A(addr[5]), .Y(n72) );
  NAND2X1 U41 ( .A(n3), .B(n72), .Y(n95) );
  NAND2X1 U43 ( .A(n12), .B(n1), .Y(n106) );
  XOR2X1 U45 ( .A(n82), .B(n2), .Y(n83) );
  NAND2X1 U46 ( .A(n1), .B(n3), .Y(n82) );
  OAI22XL U47 ( .A0(n3), .A1(n10), .B0(n70), .B1(n112), .Y(n94) );
  AOI211XL U52 ( .A0(n98), .A1(n70), .B0(n97), .C0(n104), .Y(n99) );
  OAI22XL U53 ( .A0(n96), .A1(n69), .B0(n95), .B1(n109), .Y(n97) );
  OAI22XL U54 ( .A0(n13), .A1(n72), .B0(n2), .B1(addr[1]), .Y(n98) );
  AOI221XL U55 ( .A0(n71), .A1(addr[6]), .B0(addr[5]), .B1(n94), .C0(n93), .Y(
        n96) );
  OAI21XL U58 ( .A0(addr[1]), .A1(n120), .B0(n119), .Y(n121) );
  AOI221XL U60 ( .A0(n9), .A1(n118), .B0(n93), .B1(n72), .C0(n75), .Y(n78) );
  OAI31X1 U61 ( .A0(n72), .A1(n2), .A2(n74), .B0(n73), .Y(n75) );
  OA21XL U62 ( .A0(n3), .A1(n13), .B0(n109), .Y(n74) );
  OAI21XL U63 ( .A0(n124), .A1(n85), .B0(n12), .Y(n73) );
  OAI21XL U64 ( .A0(n1), .A1(n10), .B0(n109), .Y(n110) );
  INVX4 U65 ( .A(n4), .Y(n6) );
  AOI222XL U66 ( .A0(n124), .A1(n123), .B0(n122), .B1(addr[6]), .C0(n1), .C1(
        n121), .Y(n125) );
  NOR4BBX1 U67 ( .AN(n107), .BN(n106), .C(n105), .D(n104), .Y(n127) );
  AOI222XL U68 ( .A0(n9), .A1(n90), .B0(n89), .B1(n6), .C0(n123), .C1(n69), 
        .Y(n101) );
  AOI2BB2XL U69 ( .B0(addr[5]), .B1(n92), .A0N(n120), .A1N(addr[1]), .Y(n100)
         );
  AOI32X1 U70 ( .A0(n4), .A1(n85), .A2(n9), .B0(n84), .B1(n6), .Y(n86) );
  AOI222XL U71 ( .A0(n124), .A1(n10), .B0(n83), .B1(addr[1]), .C0(n5), .C1(n13), .Y(n87) );
  OAI221X1 U72 ( .A0(n79), .A1(n72), .B0(n4), .B1(n78), .C0(n77), .Y(dout[1])
         );
  AOI32XL U73 ( .A0(addr[6]), .A1(n85), .A2(n1), .B0(n76), .B1(n72), .Y(n77)
         );
  CLKINVX3 U74 ( .A(addr[1]), .Y(n10) );
  CLKINVX3 U75 ( .A(n2), .Y(n69) );
  CLKINVX3 U76 ( .A(n3), .Y(n70) );
endmodule


module sbox2_6 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147;

  NAND2X2 U55 ( .A(n2), .B(n8), .Y(n136) );
  NAND2X2 U57 ( .A(addr[2]), .B(n16), .Y(n104) );
  NAND2X2 U60 ( .A(addr[5]), .B(addr[2]), .Y(n132) );
  NOR2X2 U61 ( .A(n13), .B(n10), .Y(n101) );
  NAND2X2 U62 ( .A(n12), .B(n82), .Y(n146) );
  NAND2X2 U63 ( .A(n3), .B(n83), .Y(n124) );
  NAND2X2 U64 ( .A(addr[6]), .B(n12), .Y(n122) );
  NAND2X2 U67 ( .A(n3), .B(n2), .Y(n133) );
  AOI222XL U1 ( .A0(n4), .A1(n14), .B0(n88), .B1(n83), .C0(n140), .C1(n10), 
        .Y(n89) );
  CLKINVX1 U2 ( .A(n121), .Y(n13) );
  OAI211X4 U3 ( .A0(n147), .A1(n146), .B0(n145), .C0(n144), .Y(dout[4]) );
  NOR2X1 U4 ( .A(n104), .B(n2), .Y(n141) );
  NOR2X1 U5 ( .A(n124), .B(n2), .Y(n140) );
  CLKBUFX4 U6 ( .A(addr[4]), .Y(n2) );
  CLKINVX1 U7 ( .A(addr[5]), .Y(n1) );
  INVX3 U8 ( .A(addr[5]), .Y(n16) );
  NAND3XL U9 ( .A(n98), .B(n97), .C(n96), .Y(dout[1]) );
  NAND2X1 U10 ( .A(addr[1]), .B(addr[6]), .Y(n121) );
  CLKINVX2 U11 ( .A(addr[1]), .Y(n12) );
  OAI221X1 U12 ( .A0(addr[1]), .A1(n136), .B0(n133), .B1(n12), .C0(n87), .Y(
        n95) );
  NAND2X4 U13 ( .A(addr[1]), .B(n82), .Y(n114) );
  INVX3 U14 ( .A(addr[6]), .Y(n82) );
  NAND2XL U15 ( .A(n102), .B(n8), .Y(n109) );
  AOI211XL U16 ( .A0(n81), .A1(n95), .B0(n94), .C0(n93), .Y(n96) );
  AOI2BB2X1 U17 ( .B0(n16), .B1(n9), .A0N(n104), .A1N(n136), .Y(n117) );
  NOR3BXL U18 ( .AN(n135), .B(n134), .C(n4), .Y(n147) );
  BUFX4 U19 ( .A(addr[3]), .Y(n3) );
  NAND2X1 U20 ( .A(n4), .B(n13), .Y(n113) );
  CLKINVX1 U21 ( .A(n146), .Y(n10) );
  CLKINVX1 U22 ( .A(n115), .Y(n4) );
  CLKINVX1 U23 ( .A(n122), .Y(n11) );
  OAI31X1 U24 ( .A0(n124), .A1(n82), .A2(n16), .B0(n123), .Y(n128) );
  OAI21XL U25 ( .A0(n16), .A1(n12), .B0(n140), .Y(n123) );
  OAI22X1 U26 ( .A0(n122), .A1(n124), .B0(n101), .B1(n132), .Y(n84) );
  INVX1 U27 ( .A(n114), .Y(n14) );
  OAI22X1 U28 ( .A0(n122), .A1(n8), .B0(n5), .B1(n121), .Y(n129) );
  NAND3X1 U29 ( .A(n5), .B(n16), .C(n12), .Y(n111) );
  NAND2X1 U30 ( .A(n8), .B(n5), .Y(n115) );
  OAI21XL U31 ( .A0(n83), .A1(n133), .B0(n135), .Y(n85) );
  OAI22XL U32 ( .A0(n117), .A1(n146), .B0(n116), .B1(n132), .Y(n118) );
  AOI222XL U33 ( .A0(n14), .A1(n115), .B0(n6), .B1(n82), .C0(n4), .C1(n10), 
        .Y(n116) );
  CLKINVX1 U34 ( .A(n104), .Y(n15) );
  OAI2BB2XL U35 ( .B0(n114), .B1(n135), .A0N(n126), .A1N(n6), .Y(n106) );
  OAI21XL U36 ( .A0(n112), .A1(n114), .B0(n111), .Y(n120) );
  OAI21XL U37 ( .A0(n133), .A1(n114), .B0(n113), .Y(n119) );
  CLKINVX1 U38 ( .A(n124), .Y(n9) );
  CLKINVX1 U39 ( .A(n136), .Y(n7) );
  CLKINVX1 U40 ( .A(n133), .Y(n6) );
  CLKINVX1 U41 ( .A(n132), .Y(n81) );
  AOI2BB1X1 U42 ( .A0N(n126), .A1N(n125), .B0(n136), .Y(n127) );
  OAI22XL U43 ( .A0(n104), .A1(n114), .B0(n101), .B1(n132), .Y(n102) );
  AO21XL U44 ( .A0(n83), .A1(n7), .B0(n141), .Y(n86) );
  AO21X1 U45 ( .A0(n8), .A1(n15), .B0(n140), .Y(n142) );
  NAND3X1 U46 ( .A(n83), .B(n5), .C(addr[5]), .Y(n135) );
  OAI22X1 U47 ( .A0(addr[5]), .A1(n121), .B0(n122), .B1(n16), .Y(n126) );
  AOI2BB1X1 U48 ( .A0N(n3), .A1N(n1), .B0(n7), .Y(n112) );
  NOR3X1 U49 ( .A(addr[1]), .B(addr[2]), .C(n16), .Y(n125) );
  AOI2BB1XL U50 ( .A0N(n92), .A1N(n91), .B0(addr[5]), .Y(n93) );
  OAI22XL U51 ( .A0(n117), .A1(n114), .B0(n89), .B1(n1), .Y(n94) );
  OAI31XL U52 ( .A0(n114), .A1(n2), .A2(n8), .B0(n90), .Y(n91) );
  OAI21XL U53 ( .A0(n6), .A1(n9), .B0(n11), .Y(n90) );
  NAND2X1 U54 ( .A(n14), .B(n2), .Y(n137) );
  OAI31XL U56 ( .A0(n101), .A1(n3), .A2(addr[2]), .B0(n113), .Y(n92) );
  OAI211X1 U58 ( .A0(n139), .A1(n16), .B0(n138), .C0(n137), .Y(n143) );
  NAND3X1 U59 ( .A(n5), .B(n16), .C(addr[6]), .Y(n138) );
  AOI2BB2X1 U65 ( .B0(n11), .B1(n8), .A0N(n12), .A1N(n136), .Y(n139) );
  OAI22XL U66 ( .A0(addr[5]), .A1(n133), .B0(n3), .B1(n132), .Y(n134) );
  OAI2BB2XL U68 ( .B0(n112), .B1(n122), .A0N(n1), .A1N(n99), .Y(n100) );
  OAI211X1 U69 ( .A0(n146), .A1(n2), .B0(n137), .C0(n113), .Y(n99) );
  NAND3X1 U70 ( .A(n11), .B(n5), .C(n3), .Y(n87) );
  AOI2BB2XL U71 ( .B0(n3), .B1(n105), .A0N(n137), .A1N(n132), .Y(n108) );
  OAI211XL U72 ( .A0(n104), .A1(n146), .B0(n103), .C0(n111), .Y(n105) );
  NAND3XL U73 ( .A(addr[5]), .B(n5), .C(n13), .Y(n103) );
  OAI22XL U74 ( .A0(n3), .A1(n114), .B0(n82), .B1(n115), .Y(n88) );
  NAND4X1 U75 ( .A(n110), .B(n109), .C(n108), .D(n107), .Y(dout[2]) );
  AOI32XL U76 ( .A0(addr[1]), .A1(addr[2]), .A2(n7), .B0(n100), .B1(n83), .Y(
        n110) );
  AOI221XL U77 ( .A0(n125), .A1(addr[4]), .B0(n141), .B1(n11), .C0(n106), .Y(
        n107) );
  AOI33XL U78 ( .A0(n11), .A1(n15), .A2(n2), .B0(n81), .B1(n146), .B2(n3), .Y(
        n145) );
  AOI222XL U79 ( .A0(n143), .A1(n83), .B0(n13), .B1(n142), .C0(n14), .C1(n141), 
        .Y(n144) );
  AOI32XL U80 ( .A0(n15), .A1(n12), .A2(n4), .B0(n10), .B1(n86), .Y(n97) );
  AOI22X1 U81 ( .A0(n13), .A1(n85), .B0(n2), .B1(n84), .Y(n98) );
  NAND2X1 U82 ( .A(n131), .B(n130), .Y(dout[3]) );
  AOI221XL U83 ( .A0(n120), .A1(n83), .B0(addr[2]), .B1(n119), .C0(n118), .Y(
        n131) );
  AOI211X1 U84 ( .A0(n15), .A1(n129), .B0(n128), .C0(n127), .Y(n130) );
  CLKINVX3 U85 ( .A(n2), .Y(n5) );
  CLKINVX3 U86 ( .A(n3), .Y(n8) );
  CLKINVX3 U87 ( .A(addr[2]), .Y(n83) );
endmodule


module sbox3_6 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134;

  NOR2X2 U35 ( .A(n8), .B(addr[3]), .Y(n109) );
  NOR2X2 U50 ( .A(addr[1]), .B(addr[6]), .Y(n108) );
  NOR2X2 U52 ( .A(n77), .B(n3), .Y(n88) );
  NOR2X2 U56 ( .A(n77), .B(n79), .Y(n95) );
  NOR2X1 U1 ( .A(n8), .B(n77), .Y(n107) );
  OAI221X1 U2 ( .A0(n125), .A1(n8), .B0(n4), .B1(addr[1]), .C0(n20), .Y(n105)
         );
  INVXL U3 ( .A(n2), .Y(n1) );
  NOR2X1 U4 ( .A(n19), .B(n4), .Y(n92) );
  NOR2X1 U5 ( .A(n10), .B(n4), .Y(n122) );
  NOR2X1 U6 ( .A(n20), .B(n4), .Y(n96) );
  CLKBUFX3 U7 ( .A(addr[2]), .Y(n4) );
  INVX1 U8 ( .A(addr[2]), .Y(n2) );
  NOR2X1 U9 ( .A(n4), .B(n3), .Y(n111) );
  BUFX4 U10 ( .A(addr[4]), .Y(n3) );
  OAI33X1 U11 ( .A0(n10), .A1(n126), .A2(n79), .B0(n8), .B1(n95), .B2(n120), 
        .Y(n80) );
  INVX3 U12 ( .A(n4), .Y(n79) );
  OAI221X1 U13 ( .A0(addr[5]), .A1(n91), .B0(n90), .B1(n5), .C0(n89), .Y(
        dout[1]) );
  NOR2X4 U14 ( .A(n78), .B(n17), .Y(n125) );
  NOR2X4 U15 ( .A(addr[3]), .B(n3), .Y(n131) );
  NOR2X4 U16 ( .A(n17), .B(addr[6]), .Y(n126) );
  INVX3 U17 ( .A(addr[1]), .Y(n17) );
  NAND2XL U18 ( .A(n95), .B(n125), .Y(n133) );
  OAI211XL U19 ( .A0(n3), .A1(n18), .B0(n129), .C0(n128), .Y(n130) );
  NAND4XL U20 ( .A(n115), .B(n114), .C(n113), .D(n112), .Y(n116) );
  CLKINVX1 U21 ( .A(n133), .Y(n15) );
  INVX1 U22 ( .A(n125), .Y(n13) );
  CLKINVX1 U23 ( .A(n107), .Y(n6) );
  NAND2X1 U24 ( .A(n19), .B(n7), .Y(n123) );
  CLKINVX1 U25 ( .A(n87), .Y(n7) );
  CLKINVX1 U26 ( .A(n121), .Y(n76) );
  CLKINVX1 U27 ( .A(n120), .Y(n14) );
  CLKINVX1 U28 ( .A(n115), .Y(n11) );
  CLKINVX1 U29 ( .A(n108), .Y(n20) );
  NOR2X1 U30 ( .A(n19), .B(n79), .Y(n104) );
  NOR2X1 U31 ( .A(n13), .B(n79), .Y(n110) );
  INVX1 U32 ( .A(n126), .Y(n16) );
  AOI21X1 U33 ( .A0(n77), .A1(n79), .B0(n95), .Y(n121) );
  OAI21XL U34 ( .A0(n111), .A1(n131), .B0(n125), .Y(n83) );
  CLKINVX1 U36 ( .A(n82), .Y(n19) );
  NOR2X1 U37 ( .A(n16), .B(n8), .Y(n87) );
  NOR2X1 U38 ( .A(n125), .B(n108), .Y(n120) );
  OAI21XL U39 ( .A0(n110), .A1(n92), .B0(n131), .Y(n101) );
  NAND2X1 U40 ( .A(n104), .B(n88), .Y(n115) );
  CLKINVX1 U41 ( .A(n88), .Y(n10) );
  CLKINVX1 U42 ( .A(n92), .Y(n18) );
  CLKINVX1 U43 ( .A(n111), .Y(n12) );
  CLKINVX1 U44 ( .A(n122), .Y(n9) );
  OR2X1 U45 ( .A(n104), .B(n96), .Y(n127) );
  OAI221X1 U46 ( .A0(n16), .A1(n12), .B0(n79), .B1(n7), .C0(n94), .Y(n99) );
  AOI221XL U47 ( .A0(n96), .A1(n3), .B0(n93), .B1(n8), .C0(n15), .Y(n94) );
  OAI21XL U48 ( .A0(n79), .A1(n20), .B0(n18), .Y(n93) );
  XNOR2X1 U49 ( .A(addr[5]), .B(addr[3]), .Y(n103) );
  CLKINVX1 U51 ( .A(addr[5]), .Y(n5) );
  OAI221X1 U53 ( .A0(n20), .A1(n12), .B0(n13), .B1(n10), .C0(n106), .Y(n117)
         );
  AOI221XL U54 ( .A0(addr[3]), .A1(n105), .B0(n104), .B1(n131), .C0(n15), .Y(
        n106) );
  CLKINVX1 U55 ( .A(addr[6]), .Y(n78) );
  NAND3X1 U57 ( .A(n4), .B(n17), .C(n109), .Y(n114) );
  NOR2X1 U58 ( .A(n78), .B(addr[1]), .Y(n82) );
  AOI32XL U59 ( .A0(n79), .A1(n77), .A2(n125), .B0(n124), .B1(n78), .Y(n129)
         );
  AOI22XL U60 ( .A0(n3), .A1(n127), .B0(n126), .B1(n131), .Y(n128) );
  OAI22XL U61 ( .A0(n3), .A1(n2), .B0(n4), .B1(n6), .Y(n124) );
  AOI222XL U62 ( .A0(n111), .A1(n126), .B0(n110), .B1(n77), .C0(n109), .C1(
        n108), .Y(n112) );
  OAI211XL U63 ( .A0(n107), .A1(n131), .B0(n2), .C0(addr[6]), .Y(n113) );
  OAI21XL U64 ( .A0(n1), .A1(addr[1]), .B0(n16), .Y(n81) );
  AOI221XL U65 ( .A0(n87), .A1(n77), .B0(n88), .B1(n126), .C0(n86), .Y(n90) );
  OAI211X1 U66 ( .A0(n85), .A1(n79), .B0(n84), .C0(n83), .Y(n86) );
  AOI222XL U67 ( .A0(n82), .A1(n77), .B0(n108), .B1(n107), .C0(n131), .C1(n17), 
        .Y(n85) );
  OAI21XL U68 ( .A0(n92), .A1(n15), .B0(addr[4]), .Y(n84) );
  AOI221XL U69 ( .A0(n126), .A1(n76), .B0(addr[3]), .B1(n127), .C0(n97), .Y(
        n98) );
  OAI22X1 U70 ( .A0(n13), .A1(n9), .B0(n6), .B1(n19), .Y(n97) );
  OAI211X1 U71 ( .A0(n20), .A1(n9), .B0(n119), .C0(n118), .Y(dout[3]) );
  AOI32XL U72 ( .A0(n126), .A1(n4), .A2(n103), .B0(n109), .B1(n110), .Y(n119)
         );
  AOI22XL U73 ( .A0(n117), .A1(n5), .B0(addr[5]), .B1(n116), .Y(n118) );
  AOI221XL U74 ( .A0(n122), .A1(n126), .B0(n96), .B1(n109), .C0(n11), .Y(n89)
         );
  AOI221XL U75 ( .A0(n131), .A1(n81), .B0(n95), .B1(n123), .C0(n80), .Y(n91)
         );
  NAND4X1 U76 ( .A(n102), .B(n114), .C(n101), .D(n100), .Y(dout[2]) );
  NAND3XL U77 ( .A(n3), .B(n125), .C(n103), .Y(n102) );
  AOI2BB2XL U78 ( .B0(addr[5]), .B1(n99), .A0N(addr[5]), .A1N(n98), .Y(n100)
         );
  OAI221X1 U79 ( .A0(n134), .A1(n5), .B0(n3), .B1(n133), .C0(n132), .Y(dout[4]) );
  AOI32XL U80 ( .A0(n131), .A1(n78), .A2(n1), .B0(n130), .B1(n5), .Y(n132) );
  AOI222XL U81 ( .A0(n76), .A1(n123), .B0(n122), .B1(addr[1]), .C0(n121), .C1(
        n14), .Y(n134) );
  CLKINVX3 U82 ( .A(n3), .Y(n8) );
  CLKINVX3 U83 ( .A(addr[3]), .Y(n77) );
endmodule


module sbox4_6 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126;

  OAI32X4 U12 ( .A0(n12), .A1(n2), .A2(addr[2]), .B0(n11), .B1(n108), .Y(n123)
         );
  OAI222X4 U20 ( .A0(addr[2]), .A1(n92), .B0(n106), .B1(n91), .C0(n90), .C1(
        n72), .Y(dout[2]) );
  OAI222X4 U33 ( .A0(addr[4]), .A1(n106), .B0(n6), .B1(n108), .C0(n2), .C1(
        n118), .Y(n83) );
  NAND2X2 U34 ( .A(addr[4]), .B(n2), .Y(n108) );
  NOR2X2 U43 ( .A(n71), .B(addr[4]), .Y(n113) );
  NOR2X2 U45 ( .A(n11), .B(n2), .Y(n111) );
  NAND2X2 U51 ( .A(n6), .B(n14), .Y(n118) );
  NOR2X2 U52 ( .A(n16), .B(addr[5]), .Y(n97) );
  NAND2X2 U53 ( .A(addr[6]), .B(addr[1]), .Y(n85) );
  NAND2X2 U54 ( .A(addr[1]), .B(n14), .Y(n116) );
  NOR2X2 U55 ( .A(n115), .B(n11), .Y(n121) );
  NAND2X2 U56 ( .A(n71), .B(n16), .Y(n115) );
  NAND2X2 U57 ( .A(addr[5]), .B(n16), .Y(n96) );
  NAND2X2 U58 ( .A(addr[6]), .B(n6), .Y(n106) );
  OAI222X1 U1 ( .A0(n12), .A1(n85), .B0(n97), .B1(n116), .C0(n16), .C1(n118), 
        .Y(n73) );
  CLKINVX1 U2 ( .A(n116), .Y(n9) );
  CLKINVX1 U3 ( .A(n71), .Y(n1) );
  CLKBUFX3 U4 ( .A(addr[3]), .Y(n2) );
  OAI31X4 U5 ( .A0(n118), .A1(n11), .A2(n16), .B0(n117), .Y(n119) );
  OAI221X1 U6 ( .A0(addr[2]), .A1(n80), .B0(n118), .B1(n105), .C0(n79), .Y(
        dout[1]) );
  INVX4 U7 ( .A(addr[5]), .Y(n11) );
  OAI31X1 U8 ( .A0(n108), .A1(addr[5]), .A2(n5), .B0(n107), .Y(n109) );
  AOI222XL U9 ( .A0(n16), .A1(n14), .B0(n113), .B1(n6), .C0(addr[1]), .C1(n71), 
        .Y(n114) );
  OAI222X1 U10 ( .A0(addr[1]), .A1(n84), .B0(n85), .B1(n74), .C0(n71), .C1(
        n107), .Y(n75) );
  NAND2XL U11 ( .A(n1), .B(addr[5]), .Y(n84) );
  AOI211XL U13 ( .A0(n83), .A1(n11), .B0(n82), .C0(n7), .Y(n92) );
  NAND2XL U14 ( .A(n16), .B(n11), .Y(n74) );
  CLKINVX1 U15 ( .A(n118), .Y(n3) );
  CLKINVX1 U16 ( .A(n115), .Y(n15) );
  CLKINVX1 U17 ( .A(n112), .Y(n4) );
  OAI21X1 U18 ( .A0(n9), .A1(n5), .B0(n72), .Y(n112) );
  AOI22X1 U19 ( .A0(n10), .A1(n111), .B0(n5), .B1(n113), .Y(n93) );
  OAI211X1 U21 ( .A0(n6), .A1(n115), .B0(n93), .C0(n8), .Y(n94) );
  CLKINVX1 U22 ( .A(n85), .Y(n10) );
  NAND2X1 U23 ( .A(n97), .B(n71), .Y(n105) );
  NAND2X1 U24 ( .A(n113), .B(n3), .Y(n98) );
  NAND2X1 U25 ( .A(n9), .B(n97), .Y(n107) );
  NAND2X1 U26 ( .A(n118), .B(n85), .Y(n110) );
  OAI21XL U27 ( .A0(n15), .A1(n11), .B0(n108), .Y(n95) );
  CLKINVX1 U28 ( .A(n84), .Y(n13) );
  CLKINVX1 U29 ( .A(addr[2]), .Y(n72) );
  OAI31X1 U30 ( .A0(n16), .A1(addr[6]), .A2(n11), .B0(n87), .Y(n88) );
  OAI21XL U31 ( .A0(n113), .A1(n12), .B0(n10), .Y(n87) );
  OAI211X1 U32 ( .A0(n76), .A1(n16), .B0(n98), .C0(n8), .Y(n77) );
  AOI222XL U35 ( .A0(addr[5]), .A1(addr[6]), .B0(n111), .B1(addr[1]), .C0(n5), 
        .C1(n2), .Y(n76) );
  NAND3XL U36 ( .A(n10), .B(n71), .C(addr[4]), .Y(n117) );
  OAI22XL U37 ( .A0(n116), .A1(n115), .B0(n1), .B1(n112), .Y(n78) );
  CLKINVX3 U38 ( .A(addr[4]), .Y(n16) );
  OAI2BB2XL U39 ( .B0(n115), .B1(n106), .A0N(n11), .A1N(n86), .Y(n89) );
  OAI221XL U40 ( .A0(n116), .A1(addr[4]), .B0(n108), .B1(addr[1]), .C0(n117), 
        .Y(n86) );
  CLKINVX1 U41 ( .A(addr[6]), .Y(n14) );
  CLKINVX1 U42 ( .A(n81), .Y(n7) );
  OAI21XL U44 ( .A0(n96), .A1(n118), .B0(n93), .Y(n82) );
  NAND3X1 U46 ( .A(n101), .B(n100), .C(n99), .Y(n102) );
  AOI32X1 U47 ( .A0(n96), .A1(n71), .A2(n9), .B0(n10), .B1(n95), .Y(n101) );
  AOI2BB2XL U48 ( .B0(n6), .B1(n121), .A0N(n98), .A1N(addr[5]), .Y(n99) );
  OAI21XL U49 ( .A0(n97), .A1(n12), .B0(n5), .Y(n100) );
  AOI2BB2XL U50 ( .B0(n5), .B1(n123), .A0N(n122), .A1N(n72), .Y(n124) );
  AOI211XL U59 ( .A0(n5), .A1(n121), .B0(n120), .C0(n119), .Y(n122) );
  OAI22XL U60 ( .A0(n116), .A1(n115), .B0(addr[5]), .B1(n114), .Y(n120) );
  CLKINVX1 U61 ( .A(n75), .Y(n8) );
  AOI32XL U62 ( .A0(n9), .A1(n96), .A2(n1), .B0(addr[1]), .B1(n121), .Y(n81)
         );
  AOI222XL U63 ( .A0(n5), .A1(n12), .B0(n121), .B1(n116), .C0(n2), .C1(n73), 
        .Y(n80) );
  AOI22XL U64 ( .A0(n78), .A1(n11), .B0(addr[2]), .B1(n77), .Y(n79) );
  NAND2XL U65 ( .A(n111), .B(addr[4]), .Y(n91) );
  AOI211X1 U66 ( .A0(n13), .A1(n110), .B0(n89), .C0(n88), .Y(n90) );
  OAI211X1 U67 ( .A0(n106), .A1(n105), .B0(n104), .C0(n103), .Y(dout[3]) );
  AOI32X1 U68 ( .A0(n2), .A1(n12), .A2(n9), .B0(n94), .B1(n72), .Y(n104) );
  AOI22XL U69 ( .A0(addr[2]), .A1(n102), .B0(n3), .B1(n123), .Y(n103) );
  OAI211X1 U70 ( .A0(addr[2]), .A1(n126), .B0(n125), .C0(n124), .Y(dout[4]) );
  AOI32X1 U71 ( .A0(n10), .A1(n12), .A2(n2), .B0(n4), .B1(n13), .Y(n125) );
  AOI221XL U72 ( .A0(n3), .A1(n111), .B0(n15), .B1(n110), .C0(n109), .Y(n126)
         );
  CLKINVX3 U73 ( .A(n106), .Y(n5) );
  CLKINVX3 U74 ( .A(addr[1]), .Y(n6) );
  CLKINVX3 U75 ( .A(n96), .Y(n12) );
  CLKINVX3 U76 ( .A(n2), .Y(n71) );
endmodule


module sbox5_6 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121;

  OAI222X4 U18 ( .A0(addr[3]), .A1(n106), .B0(n69), .B1(n90), .C0(n14), .C1(n9), .Y(n93) );
  OAI22X2 U40 ( .A0(addr[5]), .A1(n106), .B0(n70), .B1(n114), .Y(n116) );
  NOR2X2 U41 ( .A(n3), .B(addr[3]), .Y(n102) );
  NAND2X2 U45 ( .A(addr[6]), .B(n9), .Y(n114) );
  NAND2X2 U50 ( .A(n9), .B(n69), .Y(n110) );
  NAND2X2 U52 ( .A(addr[1]), .B(n69), .Y(n113) );
  NAND2X2 U54 ( .A(addr[1]), .B(addr[6]), .Y(n106) );
  NAND2X2 U55 ( .A(addr[3]), .B(n14), .Y(n121) );
  CLKINVX1 U1 ( .A(addr[5]), .Y(n1) );
  AOI221XL U2 ( .A0(n93), .A1(n1), .B0(n10), .B1(n15), .C0(n92), .Y(n105) );
  INVX3 U3 ( .A(addr[5]), .Y(n70) );
  OAI221X4 U4 ( .A0(n111), .A1(n110), .B0(n121), .B1(n114), .C0(n109), .Y(n112) );
  OAI221X4 U5 ( .A0(n14), .A1(n114), .B0(n70), .B1(n113), .C0(n120), .Y(n115)
         );
  OAI221X4 U6 ( .A0(n107), .A1(n121), .B0(n111), .B1(n113), .C0(n85), .Y(n86)
         );
  OAI31X1 U7 ( .A0(n68), .A1(addr[5]), .A2(addr[1]), .B0(n81), .Y(n73) );
  OAI32X1 U8 ( .A0(n114), .A1(addr[5]), .A2(n3), .B0(n13), .B1(n107), .Y(n79)
         );
  AOI32XL U9 ( .A0(n15), .A1(n98), .A2(n12), .B0(n2), .B1(n73), .Y(n77) );
  CLKBUFX3 U10 ( .A(addr[4]), .Y(n2) );
  CLKINVX1 U11 ( .A(n81), .Y(n5) );
  NAND2X1 U12 ( .A(n6), .B(n15), .Y(n81) );
  CLKINVX1 U13 ( .A(n110), .Y(n8) );
  CLKXOR2X2 U14 ( .A(n68), .B(n70), .Y(n94) );
  AOI2BB1X1 U15 ( .A0N(n14), .A1N(n1), .B0(n15), .Y(n111) );
  NOR2X1 U16 ( .A(n121), .B(n70), .Y(n91) );
  NOR2BX1 U17 ( .AN(n116), .B(n90), .Y(n83) );
  NAND2X1 U19 ( .A(n8), .B(n70), .Y(n120) );
  CLKINVX1 U20 ( .A(n113), .Y(n12) );
  NAND2X1 U21 ( .A(n12), .B(n70), .Y(n107) );
  CLKINVX1 U22 ( .A(n121), .Y(n13) );
  OAI31X1 U23 ( .A0(n4), .A1(n15), .A2(n113), .B0(n99), .Y(n72) );
  CLKINVX1 U24 ( .A(n106), .Y(n10) );
  OAI2BB2XL U25 ( .B0(n1), .B1(n113), .A0N(n98), .A1N(n6), .Y(n101) );
  CLKINVX1 U26 ( .A(n114), .Y(n6) );
  CLKINVX1 U27 ( .A(n90), .Y(n16) );
  CLKINVX1 U28 ( .A(addr[1]), .Y(n9) );
  CLKINVX1 U29 ( .A(addr[3]), .Y(n68) );
  CLKINVX1 U30 ( .A(addr[6]), .Y(n69) );
  AOI211X1 U31 ( .A0(n91), .A1(addr[1]), .B0(n80), .C0(n79), .Y(n89) );
  OAI2BB2XL U32 ( .B0(n111), .B1(n106), .A0N(n94), .A1N(n8), .Y(n80) );
  AOI211X1 U33 ( .A0(n102), .A1(n84), .B0(n83), .C0(n82), .Y(n85) );
  OAI21XL U34 ( .A0(n69), .A1(n1), .B0(n106), .Y(n84) );
  NOR3XL U35 ( .A(n94), .B(n3), .C(n110), .Y(n82) );
  AOI222XL U36 ( .A0(n10), .A1(n16), .B0(addr[5]), .B1(n108), .C0(n11), .C1(
        n14), .Y(n109) );
  CLKINVX1 U37 ( .A(n107), .Y(n11) );
  OAI21XL U38 ( .A0(addr[6]), .A1(addr[3]), .B0(n106), .Y(n108) );
  NAND2X1 U39 ( .A(addr[3]), .B(n3), .Y(n90) );
  NAND2X1 U42 ( .A(n2), .B(addr[5]), .Y(n98) );
  NAND2X1 U43 ( .A(n3), .B(n68), .Y(n97) );
  OAI21XL U44 ( .A0(addr[1]), .A1(n97), .B0(n96), .Y(n103) );
  AOI33XL U46 ( .A0(n3), .A1(n95), .A2(addr[5]), .B0(n94), .B1(n14), .B2(
        addr[1]), .Y(n96) );
  OAI21XL U47 ( .A0(n9), .A1(n68), .B0(n114), .Y(n95) );
  OAI21XL U48 ( .A0(addr[6]), .A1(n121), .B0(n99), .Y(n100) );
  NAND2X1 U49 ( .A(n71), .B(n8), .Y(n99) );
  XOR2X1 U51 ( .A(n4), .B(n3), .Y(n71) );
  AOI2BB2XL U53 ( .B0(n102), .B1(n116), .A0N(n2), .A1N(n75), .Y(n76) );
  AOI211X1 U56 ( .A0(n7), .A1(n3), .B0(n74), .C0(n83), .Y(n75) );
  AO22XL U57 ( .A0(n12), .A1(n13), .B0(addr[6]), .B1(n102), .Y(n74) );
  CLKINVX1 U58 ( .A(n120), .Y(n7) );
  CLKINVX1 U59 ( .A(n2), .Y(n4) );
  AO22XL U60 ( .A0(n12), .A1(n16), .B0(addr[6]), .B1(n91), .Y(n92) );
  AOI222XL U61 ( .A0(n116), .A1(n14), .B0(addr[3]), .B1(n115), .C0(n12), .C1(
        n15), .Y(n117) );
  OAI221X1 U62 ( .A0(n2), .A1(n105), .B0(n110), .B1(n121), .C0(n104), .Y(
        dout[3]) );
  AOI222XL U63 ( .A0(n2), .A1(n103), .B0(n102), .B1(n101), .C0(n100), .C1(n1), 
        .Y(n104) );
  OAI211X1 U64 ( .A0(n2), .A1(n89), .B0(n88), .C0(n87), .Y(dout[2]) );
  AOI33XL U65 ( .A0(n13), .A1(n98), .A2(n6), .B0(n3), .B1(n94), .B2(n8), .Y(
        n88) );
  AOI222XL U66 ( .A0(n5), .A1(n70), .B0(n2), .B1(n86), .C0(n91), .C1(n10), .Y(
        n87) );
  OAI211X1 U67 ( .A0(n78), .A1(n70), .B0(n77), .C0(n76), .Y(dout[1]) );
  AOI221XL U68 ( .A0(n13), .A1(addr[1]), .B0(n10), .B1(n15), .C0(n72), .Y(n78)
         );
  OAI211X1 U69 ( .A0(n121), .A1(n120), .B0(n119), .C0(n118), .Y(dout[4]) );
  AOI32XL U70 ( .A0(n15), .A1(n114), .A2(addr[5]), .B0(n2), .B1(n112), .Y(n119) );
  AOI2BB2X1 U71 ( .B0(n5), .B1(n70), .A0N(n2), .A1N(n117), .Y(n118) );
  BUFX4 U72 ( .A(addr[2]), .Y(n3) );
  CLKINVX3 U73 ( .A(n3), .Y(n14) );
  CLKINVX3 U74 ( .A(n97), .Y(n15) );
endmodule


module sbox6_6 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147;

  NAND2X2 U39 ( .A(n138), .B(addr[3]), .Y(n147) );
  NOR2X2 U47 ( .A(n15), .B(n81), .Y(n138) );
  NOR2X2 U50 ( .A(n17), .B(n4), .Y(n119) );
  NOR2X2 U58 ( .A(n11), .B(n17), .Y(n125) );
  NAND2X2 U61 ( .A(n97), .B(n103), .Y(n112) );
  NOR2X2 U62 ( .A(n85), .B(addr[1]), .Y(n103) );
  NOR2X2 U63 ( .A(n11), .B(addr[3]), .Y(n97) );
  NAND2X2 U64 ( .A(n117), .B(n131), .Y(n140) );
  NOR2X2 U65 ( .A(n5), .B(addr[3]), .Y(n131) );
  NOR2X2 U66 ( .A(n82), .B(addr[6]), .Y(n117) );
  NOR2X1 U1 ( .A(n15), .B(addr[3]), .Y(n102) );
  AOI211X1 U2 ( .A0(n7), .A1(n17), .B0(n131), .C0(n143), .Y(n121) );
  CLKINVX1 U3 ( .A(addr[3]), .Y(n1) );
  INVX3 U4 ( .A(addr[3]), .Y(n17) );
  CLKINVX1 U5 ( .A(n11), .Y(n2) );
  INVX4 U6 ( .A(n4), .Y(n11) );
  CLKBUFX3 U7 ( .A(addr[4]), .Y(n4) );
  CLKINVX1 U8 ( .A(n15), .Y(n3) );
  OAI222X1 U9 ( .A0(n91), .A1(n7), .B0(n5), .B1(n10), .C0(addr[5]), .C1(n12), 
        .Y(n92) );
  BUFX4 U10 ( .A(addr[2]), .Y(n5) );
  OAI221X1 U11 ( .A0(n85), .A1(n9), .B0(n17), .B1(n18), .C0(n86), .Y(n90) );
  INVX3 U12 ( .A(n96), .Y(n18) );
  OAI221X4 U13 ( .A0(n123), .A1(n83), .B0(n81), .B1(n7), .C0(n16), .Y(n124) );
  NOR2X4 U14 ( .A(addr[1]), .B(addr[6]), .Y(n130) );
  NOR2X4 U15 ( .A(n5), .B(addr[5]), .Y(n143) );
  INVX1 U16 ( .A(n130), .Y(n84) );
  CLKINVX1 U17 ( .A(n125), .Y(n9) );
  NAND2X1 U18 ( .A(n84), .B(n18), .Y(n105) );
  INVXL U19 ( .A(n121), .Y(n6) );
  CLKINVX1 U20 ( .A(n138), .Y(n14) );
  CLKINVX1 U21 ( .A(n117), .Y(n81) );
  CLKINVX1 U22 ( .A(n119), .Y(n12) );
  NOR2X1 U23 ( .A(n18), .B(n123), .Y(n144) );
  NOR2X1 U24 ( .A(n82), .B(n85), .Y(n96) );
  CLKINVX1 U25 ( .A(n103), .Y(n83) );
  OAI211X1 U26 ( .A0(n84), .A1(n9), .B0(n104), .C0(n112), .Y(n108) );
  OAI21XL U27 ( .A0(n103), .A1(n117), .B0(n102), .Y(n104) );
  OAI21XL U28 ( .A0(n132), .A1(n85), .B0(n1), .Y(n86) );
  AOI21X1 U29 ( .A0(n11), .A1(n102), .B0(n125), .Y(n91) );
  OAI2BB2XL U30 ( .B0(n143), .B1(n84), .A0N(n143), .A1N(n117), .Y(n118) );
  CLKINVX1 U31 ( .A(n122), .Y(n16) );
  CLKINVX1 U32 ( .A(n126), .Y(n13) );
  CLKINVX1 U33 ( .A(n97), .Y(n10) );
  NAND2BX1 U34 ( .AN(n144), .B(n137), .Y(n107) );
  CLKINVX1 U35 ( .A(addr[1]), .Y(n82) );
  NOR2X1 U36 ( .A(n18), .B(n3), .Y(n122) );
  NOR2X1 U37 ( .A(addr[1]), .B(n2), .Y(n132) );
  OAI22X1 U38 ( .A0(n12), .A1(n81), .B0(n5), .B1(n13), .Y(n88) );
  NAND2X1 U40 ( .A(n3), .B(n7), .Y(n123) );
  NAND4X1 U41 ( .A(n147), .B(n140), .C(n100), .D(n99), .Y(n101) );
  AOI222XL U42 ( .A0(n98), .A1(n15), .B0(n102), .B1(n130), .C0(n97), .C1(n105), 
        .Y(n99) );
  NAND3X1 U43 ( .A(n5), .B(n12), .C(n96), .Y(n100) );
  OAI221X1 U44 ( .A0(n17), .A1(n83), .B0(n12), .B1(n85), .C0(n13), .Y(n98) );
  AOI22X1 U45 ( .A0(n4), .A1(n115), .B0(addr[5]), .B1(n114), .Y(n129) );
  OAI21XL U46 ( .A0(n121), .A1(n84), .B0(n147), .Y(n115) );
  OAI21XL U48 ( .A0(n113), .A1(n15), .B0(n112), .Y(n114) );
  AOI221XL U49 ( .A0(n119), .A1(n82), .B0(n130), .B1(addr[3]), .C0(n111), .Y(
        n113) );
  OAI22XL U51 ( .A0(n81), .A1(n11), .B0(addr[3]), .B1(n18), .Y(n111) );
  OAI22XL U52 ( .A0(n17), .A1(n85), .B0(addr[1]), .B1(n12), .Y(n142) );
  AOI211X1 U53 ( .A0(n4), .A1(n135), .B0(n134), .C0(n133), .Y(n136) );
  OA21XL U54 ( .A0(n1), .A1(n3), .B0(n132), .Y(n133) );
  OAI2BB2XL U55 ( .B0(n2), .B1(n16), .A0N(n131), .A1N(n130), .Y(n134) );
  OAI22X1 U56 ( .A0(n5), .A1(n81), .B0(n15), .B1(n18), .Y(n135) );
  CLKINVX3 U57 ( .A(addr[5]), .Y(n7) );
  AOI2BB2X1 U59 ( .B0(n5), .B1(n130), .A0N(n3), .A1N(n83), .Y(n137) );
  NOR2X1 U60 ( .A(n83), .B(n2), .Y(n126) );
  AOI2BB2XL U67 ( .B0(n143), .B1(n90), .A0N(n89), .A1N(n7), .Y(n94) );
  AOI211X1 U68 ( .A0(n122), .A1(n4), .B0(n88), .C0(n87), .Y(n89) );
  OAI32X1 U69 ( .A0(n83), .A1(n17), .A2(n15), .B0(n14), .B1(n10), .Y(n87) );
  NAND3X1 U70 ( .A(n147), .B(n140), .C(n139), .Y(n141) );
  AOI32X1 U71 ( .A0(n5), .A1(n82), .A2(n4), .B0(n138), .B1(n11), .Y(n139) );
  AO22XL U72 ( .A0(n143), .A1(n2), .B0(n116), .B1(n11), .Y(n120) );
  OAI21XL U73 ( .A0(n3), .A1(n7), .B0(n123), .Y(n116) );
  CLKINVX1 U74 ( .A(n106), .Y(n8) );
  AOI32XL U75 ( .A0(n105), .A1(n11), .A2(n1), .B0(addr[1]), .B1(n125), .Y(n106) );
  OAI211X1 U76 ( .A0(n11), .A1(n140), .B0(n110), .C0(n109), .Y(dout[2]) );
  AOI222XL U77 ( .A0(n108), .A1(n7), .B0(n143), .B1(n8), .C0(n119), .C1(n107), 
        .Y(n109) );
  AOI2BB2XL U78 ( .B0(addr[5]), .B1(n101), .A0N(n15), .A1N(n112), .Y(n110) );
  OAI211X1 U79 ( .A0(n2), .A1(n147), .B0(n146), .C0(n145), .Y(dout[4]) );
  AOI222XL U80 ( .A0(n144), .A1(n17), .B0(n143), .B1(n142), .C0(n141), .C1(n7), 
        .Y(n145) );
  OA22X1 U81 ( .A0(n9), .A1(n137), .B0(n136), .B1(n7), .Y(n146) );
  NAND3X1 U82 ( .A(n129), .B(n128), .C(n127), .Y(dout[3]) );
  AOI32XL U83 ( .A0(n120), .A1(n17), .A2(addr[1]), .B0(n119), .B1(n118), .Y(
        n128) );
  AOI222XL U84 ( .A0(n144), .A1(n11), .B0(n126), .B1(n6), .C0(n125), .C1(n124), 
        .Y(n127) );
  NAND3BX1 U85 ( .AN(n95), .B(n94), .C(n93), .Y(dout[1]) );
  OAI222X1 U86 ( .A0(n140), .A1(n4), .B0(n112), .B1(n15), .C0(n18), .C1(n91), 
        .Y(n95) );
  AOI32XL U87 ( .A0(addr[1]), .A1(n7), .A2(n125), .B0(n130), .B1(n92), .Y(n93)
         );
  CLKINVX3 U88 ( .A(n5), .Y(n15) );
  CLKINVX3 U89 ( .A(addr[6]), .Y(n85) );
endmodule


module sbox7_6 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148;

  OAI222X4 U19 ( .A0(n20), .A1(n129), .B0(n4), .B1(n17), .C0(addr[1]), .C1(n85), .Y(n122) );
  OAI33X4 U33 ( .A0(addr[1]), .A1(n4), .A2(n5), .B0(n18), .B1(n86), .B2(n83), 
        .Y(n97) );
  NOR2X2 U44 ( .A(n84), .B(n4), .Y(n116) );
  NOR2X2 U48 ( .A(addr[1]), .B(addr[6]), .Y(n136) );
  NOR2X2 U51 ( .A(n10), .B(n84), .Y(n125) );
  NOR2X2 U52 ( .A(n18), .B(addr[3]), .Y(n131) );
  NOR2X2 U58 ( .A(n93), .B(n124), .Y(n142) );
  NOR2X2 U60 ( .A(n19), .B(addr[1]), .Y(n93) );
  NOR2X2 U62 ( .A(n87), .B(n3), .Y(n137) );
  NOR2X2 U65 ( .A(n19), .B(n21), .Y(n140) );
  NAND2X1 U1 ( .A(n3), .B(n4), .Y(n119) );
  CLKBUFX3 U2 ( .A(addr[4]), .Y(n4) );
  CLKINVX1 U3 ( .A(n87), .Y(n1) );
  CLKINVX1 U4 ( .A(n86), .Y(n2) );
  CLKBUFX3 U5 ( .A(addr[2]), .Y(n5) );
  OAI31X1 U6 ( .A0(n84), .A1(n87), .A2(n21), .B0(n117), .Y(n121) );
  NOR2X4 U7 ( .A(n21), .B(addr[6]), .Y(n124) );
  OAI22X1 U8 ( .A0(addr[1]), .A1(n85), .B0(n5), .B1(n113), .Y(n100) );
  OAI22X1 U9 ( .A0(n4), .A1(n10), .B0(addr[3]), .B1(n13), .Y(n103) );
  AOI211XL U10 ( .A0(n5), .A1(n16), .B0(n131), .C0(n130), .Y(n132) );
  NOR3XL U11 ( .A(n20), .B(addr[3]), .C(n2), .Y(n130) );
  OAI21XL U12 ( .A0(n3), .A1(n1), .B0(n119), .Y(n89) );
  BUFX4 U13 ( .A(addr[5]), .Y(n3) );
  AOI221XL U14 ( .A0(n140), .A1(n89), .B0(n109), .B1(n16), .C0(n88), .Y(n96)
         );
  CLKINVX1 U15 ( .A(n140), .Y(n18) );
  OAI2BB2XL U16 ( .B0(n142), .B1(n13), .A0N(n141), .A1N(n140), .Y(n143) );
  CLKINVX1 U17 ( .A(n125), .Y(n8) );
  CLKINVX1 U18 ( .A(n142), .Y(n16) );
  NAND2X1 U20 ( .A(n8), .B(n14), .Y(n105) );
  CLKINVX1 U21 ( .A(n123), .Y(n9) );
  CLKINVX1 U22 ( .A(n109), .Y(n12) );
  NAND2X1 U23 ( .A(n124), .B(n84), .Y(n113) );
  CLKINVX1 U24 ( .A(n137), .Y(n13) );
  NOR2X1 U25 ( .A(n13), .B(n84), .Y(n109) );
  CLKINVX1 U26 ( .A(n136), .Y(n20) );
  OAI22XL U27 ( .A0(n137), .A1(n17), .B0(n21), .B1(n12), .Y(n146) );
  OAI21X1 U28 ( .A0(n87), .A1(n8), .B0(n129), .Y(n141) );
  NAND2X1 U29 ( .A(n116), .B(n10), .Y(n129) );
  CLKINVX1 U30 ( .A(n93), .Y(n15) );
  OAI21XL U31 ( .A0(n119), .A1(n15), .B0(n118), .Y(n120) );
  OAI21XL U32 ( .A0(n125), .A1(n137), .B0(n124), .Y(n118) );
  NOR2X1 U34 ( .A(n10), .B(n85), .Y(n123) );
  CLKINVX1 U35 ( .A(n145), .Y(n85) );
  OAI22XL U36 ( .A0(n137), .A1(n113), .B0(n19), .B1(n9), .Y(n88) );
  CLKINVX1 U37 ( .A(n116), .Y(n83) );
  CLKINVX1 U38 ( .A(n131), .Y(n17) );
  CLKINVX1 U39 ( .A(n134), .Y(n14) );
  NOR2XL U40 ( .A(n125), .B(n87), .Y(n110) );
  CLKINVX1 U41 ( .A(n119), .Y(n11) );
  CLKINVX1 U42 ( .A(n103), .Y(n6) );
  OA21XL U43 ( .A0(n7), .A1(n15), .B0(n117), .Y(n102) );
  CLKINVX1 U45 ( .A(n105), .Y(n7) );
  OAI2BB1XL U46 ( .A0N(n103), .A1N(n124), .B0(n102), .Y(n104) );
  OAI22X1 U47 ( .A0(n10), .A1(n83), .B0(n4), .B1(n14), .Y(n112) );
  NOR4X1 U49 ( .A(n4), .B(addr[3]), .C(n21), .D(n86), .Y(n99) );
  XNOR2X1 U50 ( .A(addr[6]), .B(n5), .Y(n101) );
  AOI211X1 U53 ( .A0(n116), .A1(addr[6]), .B0(n115), .C0(n114), .Y(n128) );
  OAI222X1 U54 ( .A0(n111), .A1(n18), .B0(n110), .B1(n15), .C0(n20), .C1(n12), 
        .Y(n115) );
  OAI2BB2XL U55 ( .B0(n11), .B1(n113), .A0N(n21), .A1N(n112), .Y(n114) );
  OA21XL U56 ( .A0(n84), .A1(n3), .B0(n9), .Y(n111) );
  NAND2X1 U57 ( .A(n5), .B(n136), .Y(n133) );
  CLKINVX1 U59 ( .A(addr[6]), .Y(n19) );
  AOI211X1 U61 ( .A0(n131), .A1(n3), .B0(n92), .C0(n91), .Y(n95) );
  OAI221X1 U63 ( .A0(n21), .A1(n85), .B0(n18), .B1(n13), .C0(n102), .Y(n92) );
  OAI31X1 U64 ( .A0(n84), .A1(n87), .A2(n20), .B0(n90), .Y(n91) );
  AO21XL U66 ( .A0(n119), .A1(n129), .B0(addr[6]), .Y(n90) );
  NOR2X1 U67 ( .A(n87), .B(addr[3]), .Y(n145) );
  AOI21XL U68 ( .A0(addr[3]), .A1(n98), .B0(n97), .Y(n108) );
  OAI2BB1XL U69 ( .A0N(n86), .A1N(n124), .B0(n133), .Y(n98) );
  NAND3X1 U70 ( .A(n136), .B(n84), .C(n3), .Y(n117) );
  NOR2X1 U71 ( .A(addr[3]), .B(n3), .Y(n134) );
  OAI21X1 U72 ( .A0(n5), .A1(n142), .B0(n133), .Y(n138) );
  OAI22XL U73 ( .A0(n142), .A1(n83), .B0(n1), .B1(n132), .Y(n135) );
  AO21X1 U74 ( .A0(n139), .A1(n10), .B0(n138), .Y(n144) );
  OAI21XL U75 ( .A0(n2), .A1(n21), .B0(n15), .Y(n139) );
  OAI221X1 U76 ( .A0(n96), .A1(n86), .B0(n5), .B1(n95), .C0(n94), .Y(dout[1])
         );
  AOI2BB2X1 U77 ( .B0(n93), .B1(n112), .A0N(n133), .A1N(n6), .Y(n94) );
  OAI211X1 U78 ( .A0(n128), .A1(n86), .B0(n127), .C0(n126), .Y(dout[3]) );
  AOI32XL U79 ( .A0(n125), .A1(n1), .A2(n124), .B0(n123), .B1(n136), .Y(n126)
         );
  OAI31X1 U80 ( .A0(n122), .A1(n121), .A2(n120), .B0(n86), .Y(n127) );
  OAI221X1 U81 ( .A0(n3), .A1(n108), .B0(n107), .B1(n10), .C0(n106), .Y(
        dout[2]) );
  AOI32XL U82 ( .A0(n105), .A1(n86), .A2(n140), .B0(n2), .B1(n104), .Y(n106)
         );
  AOI211X1 U83 ( .A0(n101), .A1(n4), .B0(n100), .C0(n99), .Y(n107) );
  NAND2X1 U84 ( .A(n148), .B(n147), .Y(dout[4]) );
  AOI222XL U85 ( .A0(n136), .A1(n141), .B0(n3), .B1(n135), .C0(n134), .C1(n138), .Y(n148) );
  AOI222XL U86 ( .A0(n5), .A1(n146), .B0(n145), .B1(n144), .C0(n143), .C1(n86), 
        .Y(n147) );
  CLKINVX3 U87 ( .A(n3), .Y(n10) );
  CLKINVX3 U88 ( .A(addr[1]), .Y(n21) );
  CLKINVX3 U89 ( .A(addr[3]), .Y(n84) );
  CLKINVX3 U90 ( .A(n5), .Y(n86) );
  CLKINVX3 U91 ( .A(n4), .Y(n87) );
endmodule


module sbox8_6 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132;

  NAND2X2 U41 ( .A(addr[6]), .B(n6), .Y(n131) );
  NAND2X2 U48 ( .A(addr[4]), .B(n74), .Y(n123) );
  NAND2X2 U49 ( .A(n2), .B(n15), .Y(n87) );
  NAND2X2 U50 ( .A(addr[1]), .B(n16), .Y(n124) );
  NAND2X2 U54 ( .A(addr[2]), .B(n75), .Y(n116) );
  NAND2X2 U60 ( .A(addr[6]), .B(addr[1]), .Y(n105) );
  NAND2X2 U61 ( .A(n6), .B(n16), .Y(n108) );
  OAI32X1 U1 ( .A0(n16), .A1(addr[4]), .A2(n92), .B0(n115), .B1(n108), .Y(n96)
         );
  OAI31X1 U2 ( .A0(n123), .A1(addr[6]), .A2(n116), .B0(n109), .Y(n110) );
  OAI221X1 U3 ( .A0(n105), .A1(n87), .B0(addr[4]), .B1(n108), .C0(n86), .Y(n90) );
  NAND2X4 U4 ( .A(addr[4]), .B(n2), .Y(n115) );
  AOI222X1 U5 ( .A0(n88), .A1(addr[2]), .B0(n15), .B1(n10), .C0(n11), .C1(n92), 
        .Y(n114) );
  OAI222X1 U6 ( .A0(addr[2]), .A1(n126), .B0(n74), .B1(n125), .C0(n124), .C1(
        n123), .Y(n127) );
  AOI32XL U7 ( .A0(n9), .A1(n13), .A2(n2), .B0(n5), .B1(n117), .Y(n130) );
  OA21XL U8 ( .A0(n11), .A1(n75), .B0(n121), .Y(n78) );
  INVXL U9 ( .A(n119), .Y(n3) );
  INVX3 U10 ( .A(n2), .Y(n74) );
  BUFX4 U11 ( .A(addr[3]), .Y(n2) );
  CLKBUFX3 U12 ( .A(addr[5]), .Y(n1) );
  CLKINVX1 U13 ( .A(n108), .Y(n5) );
  CLKINVX1 U14 ( .A(n107), .Y(n12) );
  CLKINVX1 U15 ( .A(n93), .Y(n14) );
  NAND2X1 U16 ( .A(n74), .B(n15), .Y(n93) );
  NAND2X1 U17 ( .A(n11), .B(n75), .Y(n121) );
  OAI21XL U18 ( .A0(n115), .A1(n75), .B0(n107), .Y(n77) );
  OAI21X1 U19 ( .A0(n15), .A1(n75), .B0(n123), .Y(n88) );
  OAI31XL U20 ( .A0(n115), .A1(n6), .A2(n116), .B0(n118), .Y(n94) );
  CLKINVX1 U21 ( .A(n131), .Y(n4) );
  NAND2X1 U22 ( .A(n13), .B(n74), .Y(n107) );
  OAI22XL U23 ( .A0(n116), .A1(n123), .B0(n13), .B1(n115), .Y(n117) );
  OAI22XL U24 ( .A0(n123), .A1(n108), .B0(n131), .B1(n93), .Y(n95) );
  OAI2BB2XL U25 ( .B0(n115), .B1(n131), .A0N(n88), .A1N(n8), .Y(n89) );
  AOI211XL U26 ( .A0(n108), .A1(n105), .B0(n15), .C0(n121), .Y(n85) );
  CLKINVX1 U27 ( .A(n124), .Y(n9) );
  OAI22XL U28 ( .A0(n13), .A1(n123), .B0(n78), .B1(n87), .Y(n81) );
  NAND2BX2 U29 ( .AN(n78), .B(n74), .Y(n120) );
  NAND2XL U30 ( .A(n115), .B(n93), .Y(n104) );
  OAI2BB2XL U31 ( .B0(n106), .B1(n105), .A0N(n104), .A1N(n9), .Y(n111) );
  NOR2BXL U32 ( .AN(n123), .B(n103), .Y(n106) );
  NAND3X1 U33 ( .A(n104), .B(n6), .C(n13), .Y(n84) );
  AO21X1 U34 ( .A0(n13), .A1(n8), .B0(n101), .Y(n102) );
  OAI33X1 U35 ( .A0(n16), .A1(n74), .A2(n100), .B0(n11), .B1(n103), .B2(n124), 
        .Y(n101) );
  OA22XL U36 ( .A0(n107), .A1(n131), .B0(n120), .B1(n124), .Y(n98) );
  CLKINVX1 U37 ( .A(n125), .Y(n7) );
  OAI21XL U38 ( .A0(n9), .A1(n4), .B0(addr[4]), .Y(n86) );
  NAND2X1 U39 ( .A(n1), .B(n11), .Y(n100) );
  OAI221X1 U40 ( .A0(n124), .A1(n121), .B0(addr[1]), .B1(n120), .C0(n3), .Y(
        n128) );
  OAI31XL U42 ( .A0(n11), .A1(n6), .A2(n74), .B0(n118), .Y(n119) );
  NAND2X1 U43 ( .A(n8), .B(addr[2]), .Y(n125) );
  NAND4XL U44 ( .A(n4), .B(n1), .C(n2), .D(addr[2]), .Y(n109) );
  NAND3X1 U45 ( .A(n13), .B(n16), .C(n2), .Y(n118) );
  OAI21XL U46 ( .A0(n1), .A1(n87), .B0(n114), .Y(n76) );
  OAI22XL U47 ( .A0(n108), .A1(n120), .B0(n79), .B1(n100), .Y(n80) );
  AOI221XL U51 ( .A0(n4), .A1(n74), .B0(n8), .B1(n2), .C0(n91), .Y(n79) );
  NOR2X1 U52 ( .A(n1), .B(n2), .Y(n103) );
  NOR2X1 U53 ( .A(n87), .B(addr[6]), .Y(n91) );
  NOR2X1 U55 ( .A(n74), .B(n1), .Y(n92) );
  CLKINVX1 U56 ( .A(n100), .Y(n10) );
  OA21XL U57 ( .A0(n1), .A1(n115), .B0(n120), .Y(n132) );
  AOI221XL U58 ( .A0(n5), .A1(n2), .B0(n8), .B1(addr[4]), .C0(n122), .Y(n126)
         );
  OAI22XL U59 ( .A0(n2), .A1(n6), .B0(addr[4]), .B1(n131), .Y(n122) );
  OAI211X1 U62 ( .A0(addr[2]), .A1(n99), .B0(n98), .C0(n97), .Y(dout[2]) );
  AOI221XL U63 ( .A0(addr[2]), .A1(n96), .B0(n1), .B1(n95), .C0(n94), .Y(n97)
         );
  AOI221XL U64 ( .A0(n91), .A1(n1), .B0(n90), .B1(n75), .C0(n89), .Y(n99) );
  OAI211X1 U65 ( .A0(n132), .A1(n131), .B0(n130), .C0(n129), .Y(dout[4]) );
  AOI222XL U66 ( .A0(n128), .A1(n15), .B0(n1), .B1(n127), .C0(n12), .C1(n8), 
        .Y(n129) );
  OAI211X1 U67 ( .A0(addr[1]), .A1(n114), .B0(n113), .C0(n112), .Y(dout[3]) );
  AOI221XL U68 ( .A0(n111), .A1(n11), .B0(n12), .B1(n5), .C0(n110), .Y(n112)
         );
  AOI2BB2XL U69 ( .B0(n102), .B1(n15), .A0N(n115), .A1N(n125), .Y(n113) );
  NAND4BX1 U70 ( .AN(n85), .B(n84), .C(n83), .D(n82), .Y(dout[1]) );
  AOI221XL U71 ( .A0(n4), .A1(n81), .B0(n14), .B1(n7), .C0(n80), .Y(n82) );
  AOI22X1 U72 ( .A0(n8), .A1(n77), .B0(n9), .B1(n76), .Y(n83) );
  CLKINVX3 U73 ( .A(addr[1]), .Y(n6) );
  CLKINVX3 U74 ( .A(n105), .Y(n8) );
  CLKINVX3 U75 ( .A(addr[2]), .Y(n11) );
  CLKINVX3 U76 ( .A(n116), .Y(n13) );
  CLKINVX3 U77 ( .A(addr[4]), .Y(n15) );
  CLKINVX3 U78 ( .A(addr[6]), .Y(n16) );
  CLKINVX3 U79 ( .A(n1), .Y(n75) );
endmodule


module crp_6 ( P, R, K_sub );
  output [1:32] P;
  input [1:32] R;
  input [1:48] K_sub;
  wire   n1;
  wire   [1:48] X;

  sbox1_6 u0 ( .addr(X[1:6]), .dout({P[9], P[17], P[23], P[31]}) );
  sbox2_6 u1 ( .addr({X[7], n1, X[9:12]}), .dout({P[13], P[28], P[2], P[18]})
         );
  sbox3_6 u2 ( .addr(X[13:18]), .dout({P[24], P[16], P[30], P[6]}) );
  sbox4_6 u3 ( .addr(X[19:24]), .dout({P[26], P[20], P[10], P[1]}) );
  sbox5_6 u4 ( .addr(X[25:30]), .dout({P[8], P[14], P[25], P[3]}) );
  sbox6_6 u5 ( .addr(X[31:36]), .dout({P[4], P[29], P[11], P[19]}) );
  sbox7_6 u6 ( .addr(X[37:42]), .dout({P[32], P[12], P[22], P[7]}) );
  sbox8_6 u7 ( .addr(X[43:48]), .dout({P[5], P[27], P[15], P[21]}) );
  XOR2X1 U1 ( .A(R[1]), .B(K_sub[2]), .Y(X[2]) );
  XNOR2X1 U2 ( .A(R[5]), .B(K_sub[8]), .Y(X[8]) );
  INVX3 U3 ( .A(X[8]), .Y(n1) );
  CLKXOR2X4 U4 ( .A(R[29]), .B(K_sub[42]), .Y(X[42]) );
  CLKXOR2X4 U5 ( .A(R[16]), .B(K_sub[25]), .Y(X[25]) );
  CLKXOR2X4 U6 ( .A(R[8]), .B(K_sub[11]), .Y(X[11]) );
  CLKXOR2X4 U7 ( .A(R[22]), .B(K_sub[33]), .Y(X[33]) );
  CLKXOR2X4 U8 ( .A(R[16]), .B(K_sub[23]), .Y(X[23]) );
  CLKXOR2X4 U9 ( .A(R[10]), .B(K_sub[15]), .Y(X[15]) );
  CLKXOR2X4 U10 ( .A(R[20]), .B(K_sub[31]), .Y(X[31]) );
  CLKXOR2X4 U11 ( .A(R[31]), .B(K_sub[46]), .Y(X[46]) );
  CLKXOR2X4 U12 ( .A(R[29]), .B(K_sub[44]), .Y(X[44]) );
  CLKXOR2X4 U13 ( .A(R[12]), .B(K_sub[19]), .Y(X[19]) );
  CLKXOR2X4 U14 ( .A(R[26]), .B(K_sub[39]), .Y(X[39]) );
  CLKXOR2X4 U15 ( .A(R[20]), .B(K_sub[29]), .Y(X[29]) );
  CLKXOR2X2 U16 ( .A(R[4]), .B(K_sub[5]), .Y(X[5]) );
  CLKXOR2X2 U17 ( .A(R[15]), .B(K_sub[22]), .Y(X[22]) );
  CLKXOR2X2 U18 ( .A(R[24]), .B(K_sub[35]), .Y(X[35]) );
  CLKXOR2X2 U19 ( .A(R[21]), .B(K_sub[30]), .Y(X[30]) );
  CLKXOR2X2 U20 ( .A(R[12]), .B(K_sub[17]), .Y(X[17]) );
  CLKXOR2X2 U21 ( .A(R[32]), .B(K_sub[1]), .Y(X[1]) );
  CLKXOR2X2 U22 ( .A(R[13]), .B(K_sub[20]), .Y(X[20]) );
  CLKXOR2X2 U23 ( .A(R[18]), .B(K_sub[27]), .Y(X[27]) );
  CLKXOR2X2 U24 ( .A(R[8]), .B(K_sub[13]), .Y(X[13]) );
  CLKXOR2X2 U25 ( .A(R[5]), .B(K_sub[6]), .Y(X[6]) );
  CLKXOR2X2 U26 ( .A(R[4]), .B(K_sub[7]), .Y(X[7]) );
  CLKXOR2X2 U27 ( .A(R[24]), .B(K_sub[37]), .Y(X[37]) );
  CLKXOR2X2 U28 ( .A(R[28]), .B(K_sub[43]), .Y(X[43]) );
  CLKXOR2X2 U29 ( .A(R[1]), .B(K_sub[48]), .Y(X[48]) );
  CLKXOR2X2 U30 ( .A(R[17]), .B(K_sub[24]), .Y(X[24]) );
  CLKXOR2X2 U31 ( .A(R[9]), .B(K_sub[12]), .Y(X[12]) );
  CLKXOR2X2 U32 ( .A(R[13]), .B(K_sub[18]), .Y(X[18]) );
  CLKXOR2X2 U33 ( .A(R[25]), .B(K_sub[36]), .Y(X[36]) );
  XOR2X1 U34 ( .A(R[23]), .B(K_sub[34]), .Y(X[34]) );
  XOR2X1 U35 ( .A(R[9]), .B(K_sub[14]), .Y(X[14]) );
  XOR2X1 U36 ( .A(R[30]), .B(K_sub[45]), .Y(X[45]) );
  XOR2X1 U37 ( .A(R[21]), .B(K_sub[32]), .Y(X[32]) );
  XOR2X1 U38 ( .A(R[25]), .B(K_sub[38]), .Y(X[38]) );
  XOR2X1 U39 ( .A(R[27]), .B(K_sub[40]), .Y(X[40]) );
  XOR2X1 U40 ( .A(R[3]), .B(K_sub[4]), .Y(X[4]) );
  XOR2X1 U41 ( .A(R[11]), .B(K_sub[16]), .Y(X[16]) );
  XOR2X1 U42 ( .A(R[7]), .B(K_sub[10]), .Y(X[10]) );
  XOR2X1 U43 ( .A(R[14]), .B(K_sub[21]), .Y(X[21]) );
  XOR2X1 U44 ( .A(R[6]), .B(K_sub[9]), .Y(X[9]) );
  XOR2X1 U45 ( .A(R[2]), .B(K_sub[3]), .Y(X[3]) );
  XOR2X1 U46 ( .A(R[28]), .B(K_sub[41]), .Y(X[41]) );
  XOR2X1 U47 ( .A(R[17]), .B(K_sub[26]), .Y(X[26]) );
  XOR2X1 U48 ( .A(R[32]), .B(K_sub[47]), .Y(X[47]) );
  XOR2X1 U49 ( .A(R[19]), .B(K_sub[28]), .Y(X[28]) );
endmodule


module sbox1_5 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127;

  OAI222X4 U13 ( .A0(addr[5]), .A1(n101), .B0(n1), .B1(n100), .C0(n99), .C1(
        n72), .Y(dout[3]) );
  OAI21X2 U42 ( .A0(n4), .A1(n112), .B0(n106), .Y(n123) );
  NAND2X2 U44 ( .A(addr[6]), .B(n8), .Y(n115) );
  NAND2X2 U48 ( .A(addr[1]), .B(n13), .Y(n114) );
  OAI22X2 U49 ( .A0(n71), .A1(n12), .B0(addr[5]), .B1(n120), .Y(n85) );
  NAND2X2 U50 ( .A(n3), .B(n71), .Y(n120) );
  NOR2X2 U51 ( .A(n71), .B(n3), .Y(n124) );
  NOR2X2 U56 ( .A(n109), .B(n3), .Y(n93) );
  NAND2X2 U57 ( .A(addr[1]), .B(addr[6]), .Y(n109) );
  NAND2X2 U59 ( .A(n8), .B(n13), .Y(n112) );
  NOR2X1 U1 ( .A(n114), .B(n120), .Y(n104) );
  AOI221X4 U2 ( .A0(n7), .A1(n90), .B0(n4), .B1(n93), .C0(n102), .Y(n79) );
  NOR3X1 U3 ( .A(n2), .B(addr[6]), .C(n72), .Y(n102) );
  BUFX4 U4 ( .A(addr[4]), .Y(n2) );
  CLKBUFX3 U5 ( .A(addr[2]), .Y(n1) );
  OAI32X1 U6 ( .A0(n112), .A1(n2), .A2(n4), .B0(n115), .B1(n113), .Y(n80) );
  NOR2BXL U7 ( .AN(n118), .B(n1), .Y(n122) );
  CLKBUFX3 U8 ( .A(addr[2]), .Y(n4) );
  OAI221X4 U9 ( .A0(n88), .A1(n12), .B0(addr[5]), .B1(n87), .C0(n86), .Y(
        dout[2]) );
  OAI221X4 U10 ( .A0(addr[5]), .A1(n127), .B0(n126), .B1(n12), .C0(n125), .Y(
        dout[4]) );
  OA21XL U11 ( .A0(n95), .A1(n115), .B0(n107), .Y(n119) );
  AOI222XL U12 ( .A0(n7), .A1(n1), .B0(n2), .B1(n110), .C0(n9), .C1(n72), .Y(
        n111) );
  AOI2BB2X1 U14 ( .B0(n2), .B1(n9), .A0N(addr[4]), .A1N(n115), .Y(n91) );
  BUFX4 U15 ( .A(addr[3]), .Y(n3) );
  CLKINVX1 U16 ( .A(n112), .Y(n7) );
  CLKINVX1 U17 ( .A(n113), .Y(n69) );
  NAND2BX1 U18 ( .AN(n104), .B(n119), .Y(n84) );
  CLKXOR2X2 U19 ( .A(n70), .B(n72), .Y(n90) );
  NOR2X1 U20 ( .A(n71), .B(n70), .Y(n118) );
  OAI21XL U21 ( .A0(n70), .A1(n114), .B0(n91), .Y(n92) );
  NAND2X1 U22 ( .A(n93), .B(n71), .Y(n107) );
  NAND2X1 U23 ( .A(n72), .B(n70), .Y(n113) );
  OAI211X1 U24 ( .A0(n71), .A1(n114), .B0(n108), .C0(n107), .Y(n89) );
  CLKINVX1 U25 ( .A(n109), .Y(n9) );
  NAND2X1 U26 ( .A(n124), .B(n6), .Y(n108) );
  CLKINVX1 U27 ( .A(n114), .Y(n10) );
  CLKINVX1 U28 ( .A(n115), .Y(n6) );
  CLKINVX1 U29 ( .A(n95), .Y(n11) );
  AO22X1 U30 ( .A0(n90), .A1(n6), .B0(n70), .B1(n123), .Y(n76) );
  OAI31X1 U31 ( .A0(n72), .A1(n3), .A2(n8), .B0(n103), .Y(n105) );
  AOI31XL U32 ( .A0(n8), .A1(n72), .A2(n2), .B0(n102), .Y(n103) );
  CLKINVX1 U33 ( .A(addr[6]), .Y(n13) );
  AOI211X1 U34 ( .A0(n5), .A1(n4), .B0(n117), .C0(n116), .Y(n126) );
  CLKINVX1 U35 ( .A(n108), .Y(n5) );
  AOI211X1 U36 ( .A0(n115), .A1(n114), .B0(n113), .C0(n2), .Y(n116) );
  OAI22X1 U37 ( .A0(n120), .A1(n112), .B0(n111), .B1(n70), .Y(n117) );
  AOI211X1 U38 ( .A0(n9), .A1(n118), .B0(n81), .C0(n80), .Y(n88) );
  OAI22X1 U39 ( .A0(n91), .A1(n72), .B0(n3), .B1(n106), .Y(n81) );
  CLKINVX3 U40 ( .A(addr[5]), .Y(n12) );
  NAND2X1 U41 ( .A(n3), .B(n12), .Y(n95) );
  NAND2X1 U43 ( .A(n10), .B(n1), .Y(n106) );
  XOR2X1 U45 ( .A(n82), .B(n2), .Y(n83) );
  NAND2X1 U46 ( .A(n1), .B(n3), .Y(n82) );
  OAI22XL U47 ( .A0(n3), .A1(n8), .B0(n70), .B1(n112), .Y(n94) );
  AOI211XL U52 ( .A0(n98), .A1(n70), .B0(n97), .C0(n104), .Y(n99) );
  OAI22XL U53 ( .A0(n96), .A1(n71), .B0(n95), .B1(n109), .Y(n97) );
  OAI22XL U54 ( .A0(n13), .A1(n12), .B0(n2), .B1(addr[1]), .Y(n98) );
  AOI221XL U55 ( .A0(n11), .A1(addr[6]), .B0(addr[5]), .B1(n94), .C0(n93), .Y(
        n96) );
  OAI21XL U58 ( .A0(addr[1]), .A1(n120), .B0(n119), .Y(n121) );
  AOI221XL U60 ( .A0(n7), .A1(n118), .B0(n93), .B1(n12), .C0(n75), .Y(n78) );
  OAI31X1 U61 ( .A0(n12), .A1(n2), .A2(n74), .B0(n73), .Y(n75) );
  OA21XL U62 ( .A0(n3), .A1(n13), .B0(n109), .Y(n74) );
  OAI21XL U63 ( .A0(n124), .A1(n85), .B0(n10), .Y(n73) );
  OAI21XL U64 ( .A0(n1), .A1(n8), .B0(n109), .Y(n110) );
  INVX4 U65 ( .A(n4), .Y(n72) );
  AOI222XL U66 ( .A0(n124), .A1(n123), .B0(n122), .B1(addr[6]), .C0(n1), .C1(
        n121), .Y(n125) );
  NOR4BBX1 U67 ( .AN(n107), .BN(n106), .C(n105), .D(n104), .Y(n127) );
  AOI222XL U68 ( .A0(n7), .A1(n90), .B0(n89), .B1(n72), .C0(n123), .C1(n71), 
        .Y(n101) );
  AOI2BB2XL U69 ( .B0(addr[5]), .B1(n92), .A0N(n120), .A1N(addr[1]), .Y(n100)
         );
  AOI32X1 U70 ( .A0(n4), .A1(n85), .A2(n7), .B0(n84), .B1(n72), .Y(n86) );
  AOI222XL U71 ( .A0(n124), .A1(n8), .B0(n83), .B1(addr[1]), .C0(n69), .C1(n13), .Y(n87) );
  OAI221X1 U72 ( .A0(n79), .A1(n12), .B0(n4), .B1(n78), .C0(n77), .Y(dout[1])
         );
  AOI32XL U73 ( .A0(addr[6]), .A1(n85), .A2(n1), .B0(n76), .B1(n12), .Y(n77)
         );
  CLKINVX3 U74 ( .A(addr[1]), .Y(n8) );
  CLKINVX3 U75 ( .A(n3), .Y(n70) );
  CLKINVX3 U76 ( .A(n2), .Y(n71) );
endmodule


module sbox2_5 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147;

  NAND2X2 U55 ( .A(n2), .B(n10), .Y(n136) );
  NAND2X2 U57 ( .A(addr[2]), .B(n82), .Y(n104) );
  NAND2X2 U60 ( .A(addr[5]), .B(addr[2]), .Y(n132) );
  NOR2X2 U61 ( .A(n15), .B(n12), .Y(n101) );
  NAND2X2 U62 ( .A(n14), .B(n83), .Y(n146) );
  NAND2X2 U63 ( .A(n3), .B(n5), .Y(n124) );
  NAND2X2 U64 ( .A(addr[6]), .B(n14), .Y(n122) );
  NAND2X2 U67 ( .A(n3), .B(n2), .Y(n133) );
  AOI222XL U1 ( .A0(n9), .A1(n16), .B0(n88), .B1(n5), .C0(n140), .C1(n12), .Y(
        n89) );
  CLKINVX1 U2 ( .A(n121), .Y(n15) );
  AOI211X1 U3 ( .A0(n6), .A1(n95), .B0(n94), .C0(n93), .Y(n96) );
  NOR2X1 U4 ( .A(n104), .B(n2), .Y(n141) );
  NOR2X1 U5 ( .A(n124), .B(n2), .Y(n140) );
  CLKBUFX4 U6 ( .A(addr[4]), .Y(n2) );
  CLKINVX1 U7 ( .A(addr[5]), .Y(n1) );
  OAI22X1 U8 ( .A0(n117), .A1(n114), .B0(n89), .B1(n82), .Y(n94) );
  INVX3 U9 ( .A(addr[5]), .Y(n82) );
  OAI211X4 U10 ( .A0(n147), .A1(n146), .B0(n145), .C0(n144), .Y(dout[4]) );
  NAND2X1 U11 ( .A(addr[1]), .B(addr[6]), .Y(n121) );
  CLKINVX2 U12 ( .A(addr[1]), .Y(n14) );
  OAI221X1 U13 ( .A0(addr[1]), .A1(n136), .B0(n133), .B1(n14), .C0(n87), .Y(
        n95) );
  NAND2X4 U14 ( .A(addr[1]), .B(n83), .Y(n114) );
  INVX3 U15 ( .A(addr[6]), .Y(n83) );
  NAND2XL U16 ( .A(n102), .B(n10), .Y(n109) );
  AOI2BB2X1 U17 ( .B0(n82), .B1(n4), .A0N(n104), .A1N(n136), .Y(n117) );
  NOR3BXL U18 ( .AN(n135), .B(n134), .C(n9), .Y(n147) );
  BUFX4 U19 ( .A(addr[3]), .Y(n3) );
  NAND2X1 U20 ( .A(n9), .B(n15), .Y(n113) );
  CLKINVX1 U21 ( .A(n146), .Y(n12) );
  CLKINVX1 U22 ( .A(n115), .Y(n9) );
  CLKINVX1 U23 ( .A(n122), .Y(n13) );
  OAI31X1 U24 ( .A0(n124), .A1(n83), .A2(n82), .B0(n123), .Y(n128) );
  OAI21XL U25 ( .A0(n1), .A1(n14), .B0(n140), .Y(n123) );
  OAI22X1 U26 ( .A0(n122), .A1(n124), .B0(n101), .B1(n132), .Y(n84) );
  INVX1 U27 ( .A(n114), .Y(n16) );
  OAI22X1 U28 ( .A0(n122), .A1(n10), .B0(n81), .B1(n121), .Y(n129) );
  NAND3X1 U29 ( .A(n81), .B(n82), .C(n14), .Y(n111) );
  NAND2X1 U30 ( .A(n10), .B(n81), .Y(n115) );
  OAI21XL U31 ( .A0(n5), .A1(n133), .B0(n135), .Y(n85) );
  OAI22XL U32 ( .A0(n117), .A1(n146), .B0(n116), .B1(n132), .Y(n118) );
  AOI222XL U33 ( .A0(n16), .A1(n115), .B0(n11), .B1(n83), .C0(n9), .C1(n12), 
        .Y(n116) );
  CLKINVX1 U34 ( .A(n104), .Y(n7) );
  OAI2BB2XL U35 ( .B0(n114), .B1(n135), .A0N(n126), .A1N(n11), .Y(n106) );
  OAI21XL U36 ( .A0(n112), .A1(n114), .B0(n111), .Y(n120) );
  OAI21XL U37 ( .A0(n133), .A1(n114), .B0(n113), .Y(n119) );
  CLKINVX1 U38 ( .A(n124), .Y(n4) );
  CLKINVX1 U39 ( .A(n136), .Y(n8) );
  CLKINVX1 U40 ( .A(n133), .Y(n11) );
  CLKINVX1 U41 ( .A(n132), .Y(n6) );
  AOI2BB1X1 U42 ( .A0N(n126), .A1N(n125), .B0(n136), .Y(n127) );
  OAI22XL U43 ( .A0(n104), .A1(n114), .B0(n101), .B1(n132), .Y(n102) );
  AO21XL U44 ( .A0(n5), .A1(n8), .B0(n141), .Y(n86) );
  AO21X1 U45 ( .A0(n10), .A1(n7), .B0(n140), .Y(n142) );
  NAND3X1 U46 ( .A(n5), .B(n81), .C(addr[5]), .Y(n135) );
  OAI22X1 U47 ( .A0(addr[5]), .A1(n121), .B0(n122), .B1(n82), .Y(n126) );
  AOI2BB1X1 U48 ( .A0N(n3), .A1N(n1), .B0(n8), .Y(n112) );
  NOR3X1 U49 ( .A(addr[1]), .B(addr[2]), .C(n82), .Y(n125) );
  AOI2BB1XL U50 ( .A0N(n92), .A1N(n91), .B0(addr[5]), .Y(n93) );
  OAI31XL U51 ( .A0(n114), .A1(n2), .A2(n10), .B0(n90), .Y(n91) );
  OAI21XL U52 ( .A0(n11), .A1(n4), .B0(n13), .Y(n90) );
  NAND2X1 U53 ( .A(n16), .B(n2), .Y(n137) );
  OAI31XL U54 ( .A0(n101), .A1(n3), .A2(addr[2]), .B0(n113), .Y(n92) );
  OAI211X1 U56 ( .A0(n139), .A1(n82), .B0(n138), .C0(n137), .Y(n143) );
  NAND3X1 U58 ( .A(n81), .B(n82), .C(addr[6]), .Y(n138) );
  AOI2BB2X1 U59 ( .B0(n13), .B1(n10), .A0N(n14), .A1N(n136), .Y(n139) );
  OAI22XL U65 ( .A0(addr[5]), .A1(n133), .B0(n3), .B1(n132), .Y(n134) );
  OAI2BB2XL U66 ( .B0(n112), .B1(n122), .A0N(n1), .A1N(n99), .Y(n100) );
  OAI211X1 U68 ( .A0(n146), .A1(n2), .B0(n137), .C0(n113), .Y(n99) );
  NAND3X1 U69 ( .A(n13), .B(n81), .C(n3), .Y(n87) );
  AOI2BB2XL U70 ( .B0(n3), .B1(n105), .A0N(n137), .A1N(n132), .Y(n108) );
  OAI211XL U71 ( .A0(n104), .A1(n146), .B0(n103), .C0(n111), .Y(n105) );
  NAND3XL U72 ( .A(addr[5]), .B(n81), .C(n15), .Y(n103) );
  OAI22XL U73 ( .A0(n3), .A1(n114), .B0(n83), .B1(n115), .Y(n88) );
  NAND4X1 U74 ( .A(n110), .B(n109), .C(n108), .D(n107), .Y(dout[2]) );
  AOI32XL U75 ( .A0(addr[1]), .A1(addr[2]), .A2(n8), .B0(n100), .B1(n5), .Y(
        n110) );
  AOI221XL U76 ( .A0(n125), .A1(addr[4]), .B0(n141), .B1(n13), .C0(n106), .Y(
        n107) );
  AOI33XL U77 ( .A0(n13), .A1(n7), .A2(n2), .B0(n6), .B1(n146), .B2(n3), .Y(
        n145) );
  AOI222XL U78 ( .A0(n143), .A1(n5), .B0(n15), .B1(n142), .C0(n16), .C1(n141), 
        .Y(n144) );
  NAND3X1 U79 ( .A(n98), .B(n97), .C(n96), .Y(dout[1]) );
  AOI32XL U80 ( .A0(n7), .A1(n14), .A2(n9), .B0(n12), .B1(n86), .Y(n97) );
  AOI22X1 U81 ( .A0(n15), .A1(n85), .B0(n2), .B1(n84), .Y(n98) );
  NAND2X1 U82 ( .A(n131), .B(n130), .Y(dout[3]) );
  AOI221XL U83 ( .A0(n120), .A1(n5), .B0(addr[2]), .B1(n119), .C0(n118), .Y(
        n131) );
  AOI211X1 U84 ( .A0(n7), .A1(n129), .B0(n128), .C0(n127), .Y(n130) );
  CLKINVX3 U85 ( .A(addr[2]), .Y(n5) );
  CLKINVX3 U86 ( .A(n3), .Y(n10) );
  CLKINVX3 U87 ( .A(n2), .Y(n81) );
endmodule


module sbox3_5 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133;

  NOR2X2 U35 ( .A(n78), .B(addr[3]), .Y(n108) );
  NOR2X2 U50 ( .A(addr[1]), .B(addr[6]), .Y(n107) );
  NOR2X2 U52 ( .A(n20), .B(n2), .Y(n87) );
  NOR2X2 U56 ( .A(n20), .B(n76), .Y(n94) );
  NOR2X1 U1 ( .A(n78), .B(n20), .Y(n106) );
  OAI221X1 U2 ( .A0(n124), .A1(n78), .B0(n3), .B1(addr[1]), .C0(n13), .Y(n104)
         );
  OAI22XL U3 ( .A0(n2), .A1(n76), .B0(n3), .B1(n17), .Y(n123) );
  BUFX4 U4 ( .A(addr[4]), .Y(n2) );
  CLKBUFX3 U5 ( .A(n76), .Y(n1) );
  OAI33X1 U6 ( .A0(n19), .A1(n125), .A2(n76), .B0(n78), .B1(n94), .B2(n119), 
        .Y(n79) );
  INVX3 U7 ( .A(n3), .Y(n76) );
  NOR2X1 U8 ( .A(n12), .B(n3), .Y(n91) );
  NOR2X1 U9 ( .A(n19), .B(n3), .Y(n121) );
  NOR2X1 U10 ( .A(n13), .B(n3), .Y(n95) );
  NOR2X1 U11 ( .A(n3), .B(n2), .Y(n110) );
  CLKBUFX4 U12 ( .A(addr[2]), .Y(n3) );
  OAI221X1 U13 ( .A0(addr[5]), .A1(n90), .B0(n89), .B1(n15), .C0(n88), .Y(
        dout[1]) );
  NOR2X4 U14 ( .A(n14), .B(n9), .Y(n124) );
  NOR2X4 U15 ( .A(addr[3]), .B(n2), .Y(n130) );
  NOR2X4 U16 ( .A(n9), .B(addr[6]), .Y(n125) );
  INVX3 U17 ( .A(addr[1]), .Y(n9) );
  NAND2XL U18 ( .A(n94), .B(n124), .Y(n132) );
  OAI211XL U19 ( .A0(n2), .A1(n11), .B0(n128), .C0(n127), .Y(n129) );
  NAND4XL U20 ( .A(n114), .B(n113), .C(n112), .D(n111), .Y(n115) );
  CLKINVX1 U21 ( .A(n132), .Y(n6) );
  INVX1 U22 ( .A(n124), .Y(n4) );
  CLKINVX1 U23 ( .A(n106), .Y(n17) );
  NAND2X1 U24 ( .A(n12), .B(n7), .Y(n122) );
  CLKINVX1 U25 ( .A(n86), .Y(n7) );
  CLKINVX1 U26 ( .A(n120), .Y(n16) );
  CLKINVX1 U27 ( .A(n119), .Y(n5) );
  CLKINVX1 U28 ( .A(n114), .Y(n10) );
  CLKINVX1 U29 ( .A(n107), .Y(n13) );
  NOR2X1 U30 ( .A(n12), .B(n76), .Y(n103) );
  NOR2X1 U31 ( .A(n4), .B(n76), .Y(n109) );
  INVX1 U32 ( .A(n125), .Y(n8) );
  AOI21X1 U33 ( .A0(n20), .A1(n76), .B0(n94), .Y(n120) );
  OAI21XL U34 ( .A0(n110), .A1(n130), .B0(n124), .Y(n82) );
  CLKINVX1 U36 ( .A(n81), .Y(n12) );
  NOR2X1 U37 ( .A(n8), .B(n78), .Y(n86) );
  NOR2X1 U38 ( .A(n124), .B(n107), .Y(n119) );
  OAI21XL U39 ( .A0(n109), .A1(n91), .B0(n130), .Y(n100) );
  NAND2X1 U40 ( .A(n103), .B(n87), .Y(n114) );
  CLKINVX1 U41 ( .A(n87), .Y(n19) );
  CLKINVX1 U42 ( .A(n91), .Y(n11) );
  CLKINVX1 U43 ( .A(n110), .Y(n77) );
  CLKINVX1 U44 ( .A(n121), .Y(n18) );
  OR2X1 U45 ( .A(n103), .B(n95), .Y(n126) );
  OAI221X1 U46 ( .A0(n8), .A1(n77), .B0(n76), .B1(n7), .C0(n93), .Y(n98) );
  AOI221XL U47 ( .A0(n95), .A1(n2), .B0(n92), .B1(n78), .C0(n6), .Y(n93) );
  OAI21XL U48 ( .A0(n1), .A1(n13), .B0(n11), .Y(n92) );
  XNOR2X1 U49 ( .A(addr[5]), .B(addr[3]), .Y(n102) );
  CLKINVX1 U51 ( .A(addr[5]), .Y(n15) );
  OAI221X1 U53 ( .A0(n13), .A1(n77), .B0(n4), .B1(n19), .C0(n105), .Y(n116) );
  AOI221XL U54 ( .A0(addr[3]), .A1(n104), .B0(n103), .B1(n130), .C0(n6), .Y(
        n105) );
  CLKINVX1 U55 ( .A(addr[6]), .Y(n14) );
  NAND3X1 U57 ( .A(n3), .B(n9), .C(n108), .Y(n113) );
  NOR2X1 U58 ( .A(n14), .B(addr[1]), .Y(n81) );
  AOI32XL U59 ( .A0(n1), .A1(n20), .A2(n124), .B0(n123), .B1(n14), .Y(n128) );
  AOI22XL U60 ( .A0(n2), .A1(n126), .B0(n125), .B1(n130), .Y(n127) );
  AOI222XL U61 ( .A0(n110), .A1(n125), .B0(n109), .B1(n20), .C0(n108), .C1(
        n107), .Y(n111) );
  OAI211XL U62 ( .A0(n106), .A1(n130), .B0(n1), .C0(addr[6]), .Y(n112) );
  OAI21XL U63 ( .A0(n3), .A1(addr[1]), .B0(n8), .Y(n80) );
  AOI221XL U64 ( .A0(n86), .A1(n20), .B0(n87), .B1(n125), .C0(n85), .Y(n89) );
  OAI211X1 U65 ( .A0(n84), .A1(n76), .B0(n83), .C0(n82), .Y(n85) );
  AOI222XL U66 ( .A0(n81), .A1(n20), .B0(n107), .B1(n106), .C0(n130), .C1(n9), 
        .Y(n84) );
  OAI21XL U67 ( .A0(n91), .A1(n6), .B0(addr[4]), .Y(n83) );
  AOI221XL U68 ( .A0(n125), .A1(n16), .B0(addr[3]), .B1(n126), .C0(n96), .Y(
        n97) );
  OAI22X1 U69 ( .A0(n4), .A1(n18), .B0(n17), .B1(n12), .Y(n96) );
  OAI211X1 U70 ( .A0(n13), .A1(n18), .B0(n118), .C0(n117), .Y(dout[3]) );
  AOI32XL U71 ( .A0(n125), .A1(n3), .A2(n102), .B0(n108), .B1(n109), .Y(n118)
         );
  AOI22XL U72 ( .A0(n116), .A1(n15), .B0(addr[5]), .B1(n115), .Y(n117) );
  AOI221XL U73 ( .A0(n121), .A1(n125), .B0(n95), .B1(n108), .C0(n10), .Y(n88)
         );
  AOI221XL U74 ( .A0(n130), .A1(n80), .B0(n94), .B1(n122), .C0(n79), .Y(n90)
         );
  NAND4X1 U75 ( .A(n101), .B(n113), .C(n100), .D(n99), .Y(dout[2]) );
  NAND3XL U76 ( .A(n2), .B(n124), .C(n102), .Y(n101) );
  AOI2BB2XL U77 ( .B0(addr[5]), .B1(n98), .A0N(addr[5]), .A1N(n97), .Y(n99) );
  OAI221X1 U78 ( .A0(n133), .A1(n15), .B0(n2), .B1(n132), .C0(n131), .Y(
        dout[4]) );
  AOI32XL U79 ( .A0(n130), .A1(n14), .A2(addr[2]), .B0(n129), .B1(n15), .Y(
        n131) );
  AOI222XL U80 ( .A0(n16), .A1(n122), .B0(n121), .B1(addr[1]), .C0(n120), .C1(
        n5), .Y(n133) );
  CLKINVX3 U81 ( .A(addr[3]), .Y(n20) );
  CLKINVX3 U82 ( .A(n2), .Y(n78) );
endmodule


module sbox4_5 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126;

  OAI32X4 U12 ( .A0(n71), .A1(n2), .A2(addr[2]), .B0(n16), .B1(n108), .Y(n123)
         );
  OAI222X4 U20 ( .A0(addr[2]), .A1(n92), .B0(n106), .B1(n91), .C0(n90), .C1(
        n14), .Y(dout[2]) );
  OAI222X4 U33 ( .A0(addr[4]), .A1(n106), .B0(n6), .B1(n108), .C0(n2), .C1(
        n118), .Y(n83) );
  NAND2X2 U34 ( .A(addr[4]), .B(n2), .Y(n108) );
  NOR2X2 U43 ( .A(n12), .B(addr[4]), .Y(n113) );
  NOR2X2 U45 ( .A(n16), .B(n2), .Y(n111) );
  NAND2X2 U51 ( .A(n6), .B(n15), .Y(n118) );
  NOR2X2 U52 ( .A(n72), .B(addr[5]), .Y(n97) );
  NAND2X2 U53 ( .A(addr[6]), .B(addr[1]), .Y(n85) );
  NAND2X2 U54 ( .A(addr[1]), .B(n15), .Y(n116) );
  NOR2X2 U55 ( .A(n115), .B(n16), .Y(n121) );
  NAND2X2 U56 ( .A(n12), .B(n72), .Y(n115) );
  NAND2X2 U57 ( .A(addr[5]), .B(n72), .Y(n96) );
  NAND2X2 U58 ( .A(addr[6]), .B(n6), .Y(n106) );
  OAI222X1 U1 ( .A0(n71), .A1(n85), .B0(n97), .B1(n116), .C0(n72), .C1(n118), 
        .Y(n73) );
  CLKINVX1 U2 ( .A(n116), .Y(n9) );
  OAI31X4 U3 ( .A0(n118), .A1(n16), .A2(n72), .B0(n117), .Y(n119) );
  CLKINVX1 U4 ( .A(n12), .Y(n1) );
  CLKBUFX3 U5 ( .A(addr[3]), .Y(n2) );
  OAI221X1 U6 ( .A0(addr[2]), .A1(n80), .B0(n118), .B1(n105), .C0(n79), .Y(
        dout[1]) );
  AOI222XL U7 ( .A0(n72), .A1(n15), .B0(n113), .B1(n6), .C0(addr[1]), .C1(n12), 
        .Y(n114) );
  OAI222X1 U8 ( .A0(addr[1]), .A1(n84), .B0(n85), .B1(n74), .C0(n12), .C1(n107), .Y(n75) );
  INVX4 U9 ( .A(addr[5]), .Y(n16) );
  OAI31X1 U10 ( .A0(n108), .A1(addr[5]), .A2(n5), .B0(n107), .Y(n109) );
  NAND2XL U11 ( .A(n1), .B(addr[5]), .Y(n84) );
  AOI211XL U13 ( .A0(n83), .A1(n16), .B0(n82), .C0(n7), .Y(n92) );
  NAND2XL U14 ( .A(n72), .B(n16), .Y(n74) );
  CLKINVX1 U15 ( .A(n118), .Y(n3) );
  CLKINVX1 U16 ( .A(n115), .Y(n11) );
  CLKINVX1 U17 ( .A(n112), .Y(n4) );
  OAI21X1 U18 ( .A0(n9), .A1(n5), .B0(n14), .Y(n112) );
  AOI22X1 U19 ( .A0(n10), .A1(n111), .B0(n5), .B1(n113), .Y(n93) );
  OAI211X1 U21 ( .A0(n6), .A1(n115), .B0(n93), .C0(n8), .Y(n94) );
  CLKINVX1 U22 ( .A(n85), .Y(n10) );
  NAND2X1 U23 ( .A(n97), .B(n12), .Y(n105) );
  NAND2X1 U24 ( .A(n113), .B(n3), .Y(n98) );
  NAND2X1 U25 ( .A(n9), .B(n97), .Y(n107) );
  NAND2X1 U26 ( .A(n118), .B(n85), .Y(n110) );
  OAI21XL U27 ( .A0(n11), .A1(n16), .B0(n108), .Y(n95) );
  CLKINVX1 U28 ( .A(n84), .Y(n13) );
  CLKINVX1 U29 ( .A(addr[2]), .Y(n14) );
  OAI31X1 U30 ( .A0(n72), .A1(addr[6]), .A2(n16), .B0(n87), .Y(n88) );
  OAI21XL U31 ( .A0(n113), .A1(n71), .B0(n10), .Y(n87) );
  OAI211X1 U32 ( .A0(n76), .A1(n72), .B0(n98), .C0(n8), .Y(n77) );
  AOI222XL U35 ( .A0(addr[5]), .A1(addr[6]), .B0(n111), .B1(addr[1]), .C0(n5), 
        .C1(n2), .Y(n76) );
  NAND3XL U36 ( .A(n10), .B(n12), .C(addr[4]), .Y(n117) );
  OAI22XL U37 ( .A0(n116), .A1(n115), .B0(n1), .B1(n112), .Y(n78) );
  CLKINVX3 U38 ( .A(addr[4]), .Y(n72) );
  OAI2BB2XL U39 ( .B0(n115), .B1(n106), .A0N(n16), .A1N(n86), .Y(n89) );
  OAI221XL U40 ( .A0(n116), .A1(addr[4]), .B0(n108), .B1(addr[1]), .C0(n117), 
        .Y(n86) );
  CLKINVX1 U41 ( .A(addr[6]), .Y(n15) );
  CLKINVX1 U42 ( .A(n81), .Y(n7) );
  OAI21XL U44 ( .A0(n96), .A1(n118), .B0(n93), .Y(n82) );
  NAND3X1 U46 ( .A(n101), .B(n100), .C(n99), .Y(n102) );
  AOI32X1 U47 ( .A0(n96), .A1(n12), .A2(n9), .B0(n10), .B1(n95), .Y(n101) );
  AOI2BB2XL U48 ( .B0(n6), .B1(n121), .A0N(n98), .A1N(addr[5]), .Y(n99) );
  OAI21XL U49 ( .A0(n97), .A1(n71), .B0(n5), .Y(n100) );
  AOI2BB2XL U50 ( .B0(n5), .B1(n123), .A0N(n122), .A1N(n14), .Y(n124) );
  AOI211XL U59 ( .A0(n5), .A1(n121), .B0(n120), .C0(n119), .Y(n122) );
  OAI22XL U60 ( .A0(n116), .A1(n115), .B0(addr[5]), .B1(n114), .Y(n120) );
  CLKINVX1 U61 ( .A(n75), .Y(n8) );
  AOI32XL U62 ( .A0(n9), .A1(n96), .A2(n1), .B0(addr[1]), .B1(n121), .Y(n81)
         );
  AOI222XL U63 ( .A0(n5), .A1(n71), .B0(n121), .B1(n116), .C0(n2), .C1(n73), 
        .Y(n80) );
  AOI22XL U64 ( .A0(n78), .A1(n16), .B0(addr[2]), .B1(n77), .Y(n79) );
  NAND2XL U65 ( .A(n111), .B(addr[4]), .Y(n91) );
  AOI211X1 U66 ( .A0(n13), .A1(n110), .B0(n89), .C0(n88), .Y(n90) );
  OAI211X1 U67 ( .A0(n106), .A1(n105), .B0(n104), .C0(n103), .Y(dout[3]) );
  AOI32X1 U68 ( .A0(n2), .A1(n71), .A2(n9), .B0(n94), .B1(n14), .Y(n104) );
  AOI22XL U69 ( .A0(addr[2]), .A1(n102), .B0(n3), .B1(n123), .Y(n103) );
  OAI211X1 U70 ( .A0(addr[2]), .A1(n126), .B0(n125), .C0(n124), .Y(dout[4]) );
  AOI32X1 U71 ( .A0(n10), .A1(n71), .A2(n2), .B0(n4), .B1(n13), .Y(n125) );
  AOI221XL U72 ( .A0(n3), .A1(n111), .B0(n11), .B1(n110), .C0(n109), .Y(n126)
         );
  CLKINVX3 U73 ( .A(n106), .Y(n5) );
  CLKINVX3 U74 ( .A(addr[1]), .Y(n6) );
  CLKINVX3 U75 ( .A(n2), .Y(n12) );
  CLKINVX3 U76 ( .A(n96), .Y(n71) );
endmodule


module sbox5_5 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121;

  OAI222X4 U18 ( .A0(addr[3]), .A1(n106), .B0(n14), .B1(n90), .C0(n69), .C1(
        n68), .Y(n93) );
  OAI22X2 U40 ( .A0(addr[5]), .A1(n106), .B0(n11), .B1(n114), .Y(n116) );
  NOR2X2 U41 ( .A(n3), .B(addr[3]), .Y(n102) );
  NAND2X2 U45 ( .A(addr[6]), .B(n68), .Y(n114) );
  NAND2X2 U50 ( .A(n68), .B(n14), .Y(n110) );
  NAND2X2 U52 ( .A(addr[1]), .B(n14), .Y(n113) );
  NAND2X2 U54 ( .A(addr[1]), .B(addr[6]), .Y(n106) );
  NAND2X2 U55 ( .A(addr[3]), .B(n69), .Y(n121) );
  CLKINVX1 U1 ( .A(addr[5]), .Y(n1) );
  AOI221XL U2 ( .A0(n93), .A1(n1), .B0(n15), .B1(n5), .C0(n92), .Y(n105) );
  INVX3 U3 ( .A(addr[5]), .Y(n11) );
  OAI221X4 U4 ( .A0(n111), .A1(n110), .B0(n121), .B1(n114), .C0(n109), .Y(n112) );
  OAI221X4 U5 ( .A0(n69), .A1(n114), .B0(n11), .B1(n113), .C0(n120), .Y(n115)
         );
  OAI221X4 U6 ( .A0(n107), .A1(n121), .B0(n111), .B1(n113), .C0(n85), .Y(n86)
         );
  OAI31X1 U7 ( .A0(n6), .A1(addr[5]), .A2(addr[1]), .B0(n81), .Y(n73) );
  OAI32X1 U8 ( .A0(n114), .A1(addr[5]), .A2(n3), .B0(n7), .B1(n107), .Y(n79)
         );
  AOI32XL U9 ( .A0(n5), .A1(n98), .A2(n13), .B0(n2), .B1(n73), .Y(n77) );
  CLKBUFX3 U10 ( .A(addr[4]), .Y(n2) );
  CLKINVX1 U11 ( .A(n81), .Y(n4) );
  NAND2X1 U12 ( .A(n16), .B(n5), .Y(n81) );
  CLKINVX1 U13 ( .A(n110), .Y(n12) );
  CLKXOR2X2 U14 ( .A(n6), .B(n11), .Y(n94) );
  AOI2BB1X1 U15 ( .A0N(n69), .A1N(n1), .B0(n5), .Y(n111) );
  NOR2X1 U16 ( .A(n121), .B(n11), .Y(n91) );
  NOR2BX1 U17 ( .AN(n116), .B(n90), .Y(n83) );
  NAND2X1 U19 ( .A(n12), .B(n11), .Y(n120) );
  CLKINVX1 U20 ( .A(n113), .Y(n13) );
  NAND2X1 U21 ( .A(n13), .B(n11), .Y(n107) );
  CLKINVX1 U22 ( .A(n121), .Y(n7) );
  OAI31X1 U23 ( .A0(n70), .A1(n5), .A2(n113), .B0(n99), .Y(n72) );
  CLKINVX1 U24 ( .A(n106), .Y(n15) );
  OAI2BB2XL U25 ( .B0(n1), .B1(n113), .A0N(n98), .A1N(n16), .Y(n101) );
  CLKINVX1 U26 ( .A(n114), .Y(n16) );
  CLKINVX1 U27 ( .A(n90), .Y(n8) );
  CLKINVX1 U28 ( .A(addr[1]), .Y(n68) );
  CLKINVX1 U29 ( .A(addr[3]), .Y(n6) );
  CLKINVX1 U30 ( .A(addr[6]), .Y(n14) );
  AOI211X1 U31 ( .A0(n91), .A1(addr[1]), .B0(n80), .C0(n79), .Y(n89) );
  OAI2BB2XL U32 ( .B0(n111), .B1(n106), .A0N(n94), .A1N(n12), .Y(n80) );
  AOI211X1 U33 ( .A0(n102), .A1(n84), .B0(n83), .C0(n82), .Y(n85) );
  OAI21XL U34 ( .A0(n14), .A1(n1), .B0(n106), .Y(n84) );
  NOR3XL U35 ( .A(n94), .B(n3), .C(n110), .Y(n82) );
  AOI222XL U36 ( .A0(n15), .A1(n8), .B0(addr[5]), .B1(n108), .C0(n9), .C1(n69), 
        .Y(n109) );
  CLKINVX1 U37 ( .A(n107), .Y(n9) );
  OAI21XL U38 ( .A0(addr[6]), .A1(addr[3]), .B0(n106), .Y(n108) );
  NAND2X1 U39 ( .A(addr[3]), .B(n3), .Y(n90) );
  NAND2X1 U42 ( .A(n2), .B(addr[5]), .Y(n98) );
  NAND2X1 U43 ( .A(n3), .B(n6), .Y(n97) );
  OAI21XL U44 ( .A0(addr[1]), .A1(n97), .B0(n96), .Y(n103) );
  AOI33XL U46 ( .A0(n3), .A1(n95), .A2(addr[5]), .B0(n94), .B1(n69), .B2(
        addr[1]), .Y(n96) );
  OAI21XL U47 ( .A0(n68), .A1(n6), .B0(n114), .Y(n95) );
  OAI21XL U48 ( .A0(addr[6]), .A1(n121), .B0(n99), .Y(n100) );
  NAND2X1 U49 ( .A(n71), .B(n12), .Y(n99) );
  XOR2X1 U51 ( .A(n70), .B(n3), .Y(n71) );
  AOI2BB2XL U53 ( .B0(n102), .B1(n116), .A0N(n2), .A1N(n75), .Y(n76) );
  AOI211X1 U56 ( .A0(n10), .A1(n3), .B0(n74), .C0(n83), .Y(n75) );
  AO22XL U57 ( .A0(n13), .A1(n7), .B0(addr[6]), .B1(n102), .Y(n74) );
  CLKINVX1 U58 ( .A(n120), .Y(n10) );
  CLKINVX1 U59 ( .A(n2), .Y(n70) );
  AO22XL U60 ( .A0(n13), .A1(n8), .B0(addr[6]), .B1(n91), .Y(n92) );
  AOI222XL U61 ( .A0(n116), .A1(n69), .B0(addr[3]), .B1(n115), .C0(n13), .C1(
        n5), .Y(n117) );
  OAI221X1 U62 ( .A0(n2), .A1(n105), .B0(n110), .B1(n121), .C0(n104), .Y(
        dout[3]) );
  AOI222XL U63 ( .A0(n2), .A1(n103), .B0(n102), .B1(n101), .C0(n100), .C1(n1), 
        .Y(n104) );
  OAI211X1 U64 ( .A0(n2), .A1(n89), .B0(n88), .C0(n87), .Y(dout[2]) );
  AOI33XL U65 ( .A0(n7), .A1(n98), .A2(n16), .B0(n3), .B1(n94), .B2(n12), .Y(
        n88) );
  AOI222XL U66 ( .A0(n4), .A1(n11), .B0(n2), .B1(n86), .C0(n91), .C1(n15), .Y(
        n87) );
  OAI211X1 U67 ( .A0(n78), .A1(n11), .B0(n77), .C0(n76), .Y(dout[1]) );
  AOI221XL U68 ( .A0(n7), .A1(addr[1]), .B0(n15), .B1(n5), .C0(n72), .Y(n78)
         );
  OAI211X1 U69 ( .A0(n121), .A1(n120), .B0(n119), .C0(n118), .Y(dout[4]) );
  AOI32XL U70 ( .A0(n5), .A1(n114), .A2(addr[5]), .B0(n2), .B1(n112), .Y(n119)
         );
  AOI2BB2X1 U71 ( .B0(n4), .B1(n11), .A0N(n2), .A1N(n117), .Y(n118) );
  BUFX4 U72 ( .A(addr[2]), .Y(n3) );
  CLKINVX3 U73 ( .A(n97), .Y(n5) );
  CLKINVX3 U74 ( .A(n3), .Y(n69) );
endmodule


module sbox6_5 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147;

  NAND2X2 U39 ( .A(n138), .B(addr[3]), .Y(n147) );
  NOR2X2 U47 ( .A(n85), .B(n13), .Y(n138) );
  NOR2X2 U50 ( .A(n18), .B(n4), .Y(n119) );
  NOR2X2 U58 ( .A(n84), .B(n18), .Y(n125) );
  NAND2X2 U61 ( .A(n97), .B(n103), .Y(n112) );
  NOR2X2 U62 ( .A(n11), .B(addr[1]), .Y(n103) );
  NOR2X2 U63 ( .A(n84), .B(addr[3]), .Y(n97) );
  NAND2X2 U64 ( .A(n117), .B(n131), .Y(n140) );
  NOR2X2 U65 ( .A(n5), .B(addr[3]), .Y(n131) );
  NOR2X2 U66 ( .A(n82), .B(addr[6]), .Y(n117) );
  NOR2X1 U1 ( .A(n85), .B(addr[3]), .Y(n102) );
  OAI222X1 U2 ( .A0(n91), .A1(n83), .B0(n2), .B1(n81), .C0(addr[5]), .C1(n16), 
        .Y(n92) );
  CLKINVX1 U3 ( .A(n84), .Y(n1) );
  INVX4 U4 ( .A(n4), .Y(n84) );
  CLKBUFX3 U5 ( .A(addr[4]), .Y(n4) );
  CLKINVX1 U6 ( .A(n85), .Y(n2) );
  BUFX4 U7 ( .A(addr[2]), .Y(n5) );
  CLKINVX1 U8 ( .A(addr[3]), .Y(n3) );
  OAI22X1 U9 ( .A0(n18), .A1(n11), .B0(addr[1]), .B1(n16), .Y(n142) );
  AOI211X1 U10 ( .A0(n83), .A1(n18), .B0(n131), .C0(n143), .Y(n121) );
  INVX3 U11 ( .A(addr[3]), .Y(n18) );
  OAI221X1 U12 ( .A0(n11), .A1(n17), .B0(n18), .B1(n8), .C0(n86), .Y(n90) );
  INVX3 U13 ( .A(n96), .Y(n8) );
  OAI221X4 U14 ( .A0(n123), .A1(n10), .B0(n13), .B1(n83), .C0(n7), .Y(n124) );
  NOR2X4 U15 ( .A(addr[1]), .B(addr[6]), .Y(n130) );
  NOR2X4 U16 ( .A(n5), .B(addr[5]), .Y(n143) );
  INVX1 U17 ( .A(n130), .Y(n14) );
  CLKINVX1 U18 ( .A(n125), .Y(n17) );
  NAND2X1 U19 ( .A(n14), .B(n8), .Y(n105) );
  INVXL U20 ( .A(n121), .Y(n15) );
  CLKINVX1 U21 ( .A(n138), .Y(n12) );
  CLKINVX1 U22 ( .A(n117), .Y(n13) );
  CLKINVX1 U23 ( .A(n119), .Y(n16) );
  NOR2X1 U24 ( .A(n8), .B(n123), .Y(n144) );
  NOR2X1 U25 ( .A(n82), .B(n11), .Y(n96) );
  CLKINVX1 U26 ( .A(n103), .Y(n10) );
  OAI211X1 U27 ( .A0(n14), .A1(n17), .B0(n104), .C0(n112), .Y(n108) );
  OAI21XL U28 ( .A0(n103), .A1(n117), .B0(n102), .Y(n104) );
  OAI21XL U29 ( .A0(n132), .A1(n11), .B0(n3), .Y(n86) );
  AOI21X1 U30 ( .A0(n84), .A1(n102), .B0(n125), .Y(n91) );
  OAI2BB2XL U31 ( .B0(n143), .B1(n14), .A0N(n143), .A1N(n117), .Y(n118) );
  CLKINVX1 U32 ( .A(n122), .Y(n7) );
  CLKINVX1 U33 ( .A(n126), .Y(n9) );
  CLKINVX1 U34 ( .A(n97), .Y(n81) );
  NAND2BX1 U35 ( .AN(n144), .B(n137), .Y(n107) );
  CLKINVX1 U36 ( .A(addr[1]), .Y(n82) );
  NOR2X1 U37 ( .A(n8), .B(n2), .Y(n122) );
  NOR2X1 U38 ( .A(addr[1]), .B(n1), .Y(n132) );
  OAI22X1 U40 ( .A0(n16), .A1(n13), .B0(n5), .B1(n9), .Y(n88) );
  NAND2X1 U41 ( .A(n5), .B(n83), .Y(n123) );
  NAND4X1 U42 ( .A(n147), .B(n140), .C(n100), .D(n99), .Y(n101) );
  AOI222XL U43 ( .A0(n98), .A1(n85), .B0(n102), .B1(n130), .C0(n97), .C1(n105), 
        .Y(n99) );
  NAND3X1 U44 ( .A(n5), .B(n16), .C(n96), .Y(n100) );
  OAI221X1 U45 ( .A0(n18), .A1(n10), .B0(n16), .B1(n11), .C0(n9), .Y(n98) );
  AOI22X1 U46 ( .A0(n4), .A1(n115), .B0(addr[5]), .B1(n114), .Y(n129) );
  OAI21XL U48 ( .A0(n121), .A1(n14), .B0(n147), .Y(n115) );
  OAI21XL U49 ( .A0(n113), .A1(n85), .B0(n112), .Y(n114) );
  AOI221XL U51 ( .A0(n119), .A1(n82), .B0(n130), .B1(addr[3]), .C0(n111), .Y(
        n113) );
  OAI22XL U52 ( .A0(n13), .A1(n84), .B0(addr[3]), .B1(n8), .Y(n111) );
  AOI211X1 U53 ( .A0(n4), .A1(n135), .B0(n134), .C0(n133), .Y(n136) );
  OA21XL U54 ( .A0(n3), .A1(n2), .B0(n132), .Y(n133) );
  OAI2BB2XL U55 ( .B0(n1), .B1(n7), .A0N(n131), .A1N(n130), .Y(n134) );
  OAI22X1 U56 ( .A0(n5), .A1(n13), .B0(n85), .B1(n8), .Y(n135) );
  CLKINVX3 U57 ( .A(addr[5]), .Y(n83) );
  AOI2BB2X1 U59 ( .B0(n5), .B1(n130), .A0N(n2), .A1N(n10), .Y(n137) );
  NOR2X1 U60 ( .A(n10), .B(n1), .Y(n126) );
  AOI2BB2XL U67 ( .B0(n143), .B1(n90), .A0N(n89), .A1N(n83), .Y(n94) );
  AOI211X1 U68 ( .A0(n122), .A1(n4), .B0(n88), .C0(n87), .Y(n89) );
  OAI32X1 U69 ( .A0(n10), .A1(n18), .A2(n85), .B0(n12), .B1(n81), .Y(n87) );
  NAND3X1 U70 ( .A(n147), .B(n140), .C(n139), .Y(n141) );
  AOI32X1 U71 ( .A0(n5), .A1(n82), .A2(n4), .B0(n138), .B1(n84), .Y(n139) );
  AO22XL U72 ( .A0(n143), .A1(n1), .B0(n116), .B1(n84), .Y(n120) );
  OAI21XL U73 ( .A0(n2), .A1(n83), .B0(n123), .Y(n116) );
  CLKINVX1 U74 ( .A(n106), .Y(n6) );
  AOI32XL U75 ( .A0(n105), .A1(n84), .A2(n3), .B0(addr[1]), .B1(n125), .Y(n106) );
  OAI211X1 U76 ( .A0(n84), .A1(n140), .B0(n110), .C0(n109), .Y(dout[2]) );
  AOI222XL U77 ( .A0(n108), .A1(n83), .B0(n143), .B1(n6), .C0(n119), .C1(n107), 
        .Y(n109) );
  AOI2BB2XL U78 ( .B0(addr[5]), .B1(n101), .A0N(n85), .A1N(n112), .Y(n110) );
  OAI211X1 U79 ( .A0(n1), .A1(n147), .B0(n146), .C0(n145), .Y(dout[4]) );
  AOI222XL U80 ( .A0(n144), .A1(n18), .B0(n143), .B1(n142), .C0(n141), .C1(n83), .Y(n145) );
  OA22X1 U81 ( .A0(n17), .A1(n137), .B0(n136), .B1(n83), .Y(n146) );
  NAND3X1 U82 ( .A(n129), .B(n128), .C(n127), .Y(dout[3]) );
  AOI32XL U83 ( .A0(n120), .A1(n18), .A2(addr[1]), .B0(n119), .B1(n118), .Y(
        n128) );
  AOI222XL U84 ( .A0(n144), .A1(n84), .B0(n126), .B1(n15), .C0(n125), .C1(n124), .Y(n127) );
  NAND3BX1 U85 ( .AN(n95), .B(n94), .C(n93), .Y(dout[1]) );
  OAI222X1 U86 ( .A0(n140), .A1(n4), .B0(n112), .B1(n85), .C0(n8), .C1(n91), 
        .Y(n95) );
  AOI32XL U87 ( .A0(addr[1]), .A1(n83), .A2(n125), .B0(n130), .B1(n92), .Y(n93) );
  CLKINVX3 U88 ( .A(addr[6]), .Y(n11) );
  CLKINVX3 U89 ( .A(n5), .Y(n85) );
endmodule


module sbox7_5 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148;

  OAI222X4 U19 ( .A0(n11), .A1(n129), .B0(n4), .B1(n7), .C0(addr[1]), .C1(n13), 
        .Y(n122) );
  OAI33X4 U33 ( .A0(addr[1]), .A1(n4), .A2(n5), .B0(n8), .B1(n85), .B2(n19), 
        .Y(n97) );
  NOR2X2 U44 ( .A(n87), .B(n4), .Y(n116) );
  NOR2X2 U48 ( .A(addr[1]), .B(addr[6]), .Y(n136) );
  NOR2X2 U51 ( .A(n83), .B(n87), .Y(n125) );
  NOR2X2 U52 ( .A(n8), .B(addr[3]), .Y(n131) );
  NOR2X2 U58 ( .A(n93), .B(n124), .Y(n142) );
  NOR2X2 U60 ( .A(n86), .B(addr[1]), .Y(n93) );
  NOR2X2 U62 ( .A(n17), .B(n3), .Y(n137) );
  NOR2X2 U65 ( .A(n86), .B(n9), .Y(n140) );
  NAND2X1 U1 ( .A(n3), .B(n4), .Y(n119) );
  CLKBUFX3 U2 ( .A(addr[4]), .Y(n4) );
  CLKINVX1 U3 ( .A(n17), .Y(n1) );
  CLKINVX1 U4 ( .A(n85), .Y(n2) );
  CLKBUFX3 U5 ( .A(addr[2]), .Y(n5) );
  OAI31X1 U6 ( .A0(n87), .A1(n17), .A2(n9), .B0(n117), .Y(n121) );
  NOR2X4 U7 ( .A(n9), .B(addr[6]), .Y(n124) );
  OAI22X1 U8 ( .A0(addr[1]), .A1(n13), .B0(n5), .B1(n113), .Y(n100) );
  OAI22X1 U9 ( .A0(n4), .A1(n83), .B0(addr[3]), .B1(n16), .Y(n103) );
  AOI211XL U10 ( .A0(n5), .A1(n6), .B0(n131), .C0(n130), .Y(n132) );
  NOR3XL U11 ( .A(n11), .B(addr[3]), .C(n2), .Y(n130) );
  OAI21XL U12 ( .A0(n3), .A1(n1), .B0(n119), .Y(n89) );
  BUFX4 U13 ( .A(addr[5]), .Y(n3) );
  AOI221XL U14 ( .A0(n140), .A1(n89), .B0(n109), .B1(n6), .C0(n88), .Y(n96) );
  CLKINVX1 U15 ( .A(n140), .Y(n8) );
  OAI2BB2XL U16 ( .B0(n142), .B1(n16), .A0N(n141), .A1N(n140), .Y(n143) );
  CLKINVX1 U17 ( .A(n125), .Y(n21) );
  CLKINVX1 U18 ( .A(n142), .Y(n6) );
  NAND2X1 U20 ( .A(n21), .B(n84), .Y(n105) );
  CLKINVX1 U21 ( .A(n123), .Y(n12) );
  CLKINVX1 U22 ( .A(n109), .Y(n15) );
  NAND2X1 U23 ( .A(n124), .B(n87), .Y(n113) );
  CLKINVX1 U24 ( .A(n137), .Y(n16) );
  NOR2X1 U25 ( .A(n16), .B(n87), .Y(n109) );
  CLKINVX1 U26 ( .A(n136), .Y(n11) );
  OAI22XL U27 ( .A0(n137), .A1(n7), .B0(n9), .B1(n15), .Y(n146) );
  OAI21X1 U28 ( .A0(n17), .A1(n21), .B0(n129), .Y(n141) );
  NAND2X1 U29 ( .A(n116), .B(n83), .Y(n129) );
  CLKINVX1 U30 ( .A(n93), .Y(n10) );
  OAI21XL U31 ( .A0(n119), .A1(n10), .B0(n118), .Y(n120) );
  OAI21XL U32 ( .A0(n125), .A1(n137), .B0(n124), .Y(n118) );
  NOR2X1 U34 ( .A(n83), .B(n13), .Y(n123) );
  CLKINVX1 U35 ( .A(n145), .Y(n13) );
  OAI22XL U36 ( .A0(n137), .A1(n113), .B0(n86), .B1(n12), .Y(n88) );
  CLKINVX1 U37 ( .A(n116), .Y(n19) );
  CLKINVX1 U38 ( .A(n131), .Y(n7) );
  CLKINVX1 U39 ( .A(n134), .Y(n84) );
  NOR2XL U40 ( .A(n125), .B(n17), .Y(n110) );
  CLKINVX1 U41 ( .A(n119), .Y(n18) );
  CLKINVX1 U42 ( .A(n103), .Y(n14) );
  OA21XL U43 ( .A0(n20), .A1(n10), .B0(n117), .Y(n102) );
  CLKINVX1 U45 ( .A(n105), .Y(n20) );
  OAI2BB1XL U46 ( .A0N(n103), .A1N(n124), .B0(n102), .Y(n104) );
  OAI22X1 U47 ( .A0(n83), .A1(n19), .B0(n4), .B1(n84), .Y(n112) );
  NOR4X1 U49 ( .A(n4), .B(addr[3]), .C(n9), .D(n85), .Y(n99) );
  XNOR2X1 U50 ( .A(addr[6]), .B(n5), .Y(n101) );
  AOI211X1 U53 ( .A0(n116), .A1(addr[6]), .B0(n115), .C0(n114), .Y(n128) );
  OAI222X1 U54 ( .A0(n111), .A1(n8), .B0(n110), .B1(n10), .C0(n11), .C1(n15), 
        .Y(n115) );
  OAI2BB2XL U55 ( .B0(n18), .B1(n113), .A0N(n9), .A1N(n112), .Y(n114) );
  OA21XL U56 ( .A0(n87), .A1(n3), .B0(n12), .Y(n111) );
  NAND2X1 U57 ( .A(n5), .B(n136), .Y(n133) );
  CLKINVX1 U59 ( .A(addr[6]), .Y(n86) );
  AOI211X1 U61 ( .A0(n131), .A1(n3), .B0(n92), .C0(n91), .Y(n95) );
  OAI221X1 U63 ( .A0(n9), .A1(n13), .B0(n8), .B1(n16), .C0(n102), .Y(n92) );
  OAI31X1 U64 ( .A0(n87), .A1(n17), .A2(n11), .B0(n90), .Y(n91) );
  AO21XL U66 ( .A0(n119), .A1(n129), .B0(addr[6]), .Y(n90) );
  NOR2X1 U67 ( .A(n17), .B(addr[3]), .Y(n145) );
  AOI21XL U68 ( .A0(addr[3]), .A1(n98), .B0(n97), .Y(n108) );
  OAI2BB1XL U69 ( .A0N(n85), .A1N(n124), .B0(n133), .Y(n98) );
  NAND3X1 U70 ( .A(n136), .B(n87), .C(n3), .Y(n117) );
  NOR2X1 U71 ( .A(addr[3]), .B(n3), .Y(n134) );
  OAI21X1 U72 ( .A0(n5), .A1(n142), .B0(n133), .Y(n138) );
  OAI22XL U73 ( .A0(n142), .A1(n19), .B0(n1), .B1(n132), .Y(n135) );
  AO21X1 U74 ( .A0(n139), .A1(n83), .B0(n138), .Y(n144) );
  OAI21XL U75 ( .A0(n2), .A1(n9), .B0(n10), .Y(n139) );
  OAI221X1 U76 ( .A0(n96), .A1(n85), .B0(n5), .B1(n95), .C0(n94), .Y(dout[1])
         );
  AOI2BB2X1 U77 ( .B0(n93), .B1(n112), .A0N(n133), .A1N(n14), .Y(n94) );
  OAI211X1 U78 ( .A0(n128), .A1(n85), .B0(n127), .C0(n126), .Y(dout[3]) );
  AOI32XL U79 ( .A0(n125), .A1(n1), .A2(n124), .B0(n123), .B1(n136), .Y(n126)
         );
  OAI31X1 U80 ( .A0(n122), .A1(n121), .A2(n120), .B0(n85), .Y(n127) );
  OAI221X1 U81 ( .A0(n3), .A1(n108), .B0(n107), .B1(n83), .C0(n106), .Y(
        dout[2]) );
  AOI32XL U82 ( .A0(n105), .A1(n85), .A2(n140), .B0(n2), .B1(n104), .Y(n106)
         );
  AOI211X1 U83 ( .A0(n101), .A1(n4), .B0(n100), .C0(n99), .Y(n107) );
  NAND2X1 U84 ( .A(n148), .B(n147), .Y(dout[4]) );
  AOI222XL U85 ( .A0(n136), .A1(n141), .B0(n3), .B1(n135), .C0(n134), .C1(n138), .Y(n148) );
  AOI222XL U86 ( .A0(n5), .A1(n146), .B0(n145), .B1(n144), .C0(n143), .C1(n85), 
        .Y(n147) );
  CLKINVX3 U87 ( .A(addr[1]), .Y(n9) );
  CLKINVX3 U88 ( .A(n4), .Y(n17) );
  CLKINVX3 U89 ( .A(n3), .Y(n83) );
  CLKINVX3 U90 ( .A(n5), .Y(n85) );
  CLKINVX3 U91 ( .A(addr[3]), .Y(n87) );
endmodule


module sbox8_5 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132;

  NAND2X2 U41 ( .A(addr[6]), .B(n14), .Y(n131) );
  NAND2X2 U48 ( .A(addr[4]), .B(n7), .Y(n123) );
  NAND2X2 U49 ( .A(n2), .B(n4), .Y(n87) );
  NAND2X2 U50 ( .A(addr[1]), .B(n75), .Y(n124) );
  NAND2X2 U54 ( .A(addr[2]), .B(n74), .Y(n116) );
  NAND2X2 U60 ( .A(addr[6]), .B(addr[1]), .Y(n105) );
  NAND2X2 U61 ( .A(n14), .B(n75), .Y(n108) );
  OAI31X1 U1 ( .A0(n123), .A1(addr[6]), .A2(n116), .B0(n109), .Y(n110) );
  AOI222X1 U2 ( .A0(n88), .A1(addr[2]), .B0(n4), .B1(n8), .C0(n9), .C1(n92), 
        .Y(n114) );
  OAI222X1 U3 ( .A0(addr[2]), .A1(n126), .B0(n7), .B1(n125), .C0(n124), .C1(
        n123), .Y(n127) );
  NAND2X4 U4 ( .A(addr[4]), .B(n2), .Y(n115) );
  OAI32X1 U5 ( .A0(n75), .A1(addr[4]), .A2(n92), .B0(n115), .B1(n108), .Y(n96)
         );
  OAI221X1 U6 ( .A0(n105), .A1(n87), .B0(addr[4]), .B1(n108), .C0(n86), .Y(n90) );
  AOI32XL U7 ( .A0(n16), .A1(n10), .A2(n2), .B0(n13), .B1(n117), .Y(n130) );
  OA21XL U8 ( .A0(n9), .A1(n74), .B0(n121), .Y(n78) );
  INVXL U9 ( .A(n119), .Y(n5) );
  INVX3 U10 ( .A(n2), .Y(n7) );
  BUFX4 U11 ( .A(addr[3]), .Y(n2) );
  CLKBUFX3 U12 ( .A(addr[5]), .Y(n1) );
  CLKINVX1 U13 ( .A(n108), .Y(n13) );
  CLKINVX1 U14 ( .A(n107), .Y(n6) );
  CLKINVX1 U15 ( .A(n93), .Y(n3) );
  NAND2X1 U16 ( .A(n7), .B(n4), .Y(n93) );
  NAND2X1 U17 ( .A(n9), .B(n74), .Y(n121) );
  OAI21XL U18 ( .A0(n115), .A1(n74), .B0(n107), .Y(n77) );
  OAI21X1 U19 ( .A0(n4), .A1(n74), .B0(n123), .Y(n88) );
  OAI31XL U20 ( .A0(n115), .A1(n14), .A2(n116), .B0(n118), .Y(n94) );
  CLKINVX1 U21 ( .A(n131), .Y(n12) );
  NAND2X1 U22 ( .A(n10), .B(n7), .Y(n107) );
  OAI22XL U23 ( .A0(n116), .A1(n123), .B0(n10), .B1(n115), .Y(n117) );
  OAI22XL U24 ( .A0(n123), .A1(n108), .B0(n131), .B1(n93), .Y(n95) );
  OAI2BB2XL U25 ( .B0(n115), .B1(n131), .A0N(n88), .A1N(n15), .Y(n89) );
  AOI211XL U26 ( .A0(n108), .A1(n105), .B0(n4), .C0(n121), .Y(n85) );
  CLKINVX1 U27 ( .A(n124), .Y(n16) );
  OAI22XL U28 ( .A0(n10), .A1(n123), .B0(n78), .B1(n87), .Y(n81) );
  NAND2BX2 U29 ( .AN(n78), .B(n7), .Y(n120) );
  NAND2XL U30 ( .A(n115), .B(n93), .Y(n104) );
  OAI2BB2XL U31 ( .B0(n106), .B1(n105), .A0N(n104), .A1N(n16), .Y(n111) );
  NOR2BXL U32 ( .AN(n123), .B(n103), .Y(n106) );
  NAND3X1 U33 ( .A(n104), .B(n14), .C(n10), .Y(n84) );
  AO21X1 U34 ( .A0(n10), .A1(n15), .B0(n101), .Y(n102) );
  OAI33X1 U35 ( .A0(n75), .A1(n7), .A2(n100), .B0(n9), .B1(n103), .B2(n124), 
        .Y(n101) );
  OA22XL U36 ( .A0(n107), .A1(n131), .B0(n120), .B1(n124), .Y(n98) );
  CLKINVX1 U37 ( .A(n125), .Y(n11) );
  OAI21XL U38 ( .A0(n16), .A1(n12), .B0(addr[4]), .Y(n86) );
  NAND2X1 U39 ( .A(n1), .B(n9), .Y(n100) );
  OAI221X1 U40 ( .A0(n124), .A1(n121), .B0(addr[1]), .B1(n120), .C0(n5), .Y(
        n128) );
  OAI31XL U42 ( .A0(n9), .A1(n14), .A2(n7), .B0(n118), .Y(n119) );
  NAND2X1 U43 ( .A(n15), .B(addr[2]), .Y(n125) );
  NAND4XL U44 ( .A(n12), .B(n1), .C(n2), .D(addr[2]), .Y(n109) );
  NAND3X1 U45 ( .A(n10), .B(n75), .C(n2), .Y(n118) );
  OAI21XL U46 ( .A0(n1), .A1(n87), .B0(n114), .Y(n76) );
  OAI22XL U47 ( .A0(n108), .A1(n120), .B0(n79), .B1(n100), .Y(n80) );
  AOI221XL U51 ( .A0(n12), .A1(n7), .B0(n15), .B1(n2), .C0(n91), .Y(n79) );
  NOR2X1 U52 ( .A(n1), .B(n2), .Y(n103) );
  NOR2X1 U53 ( .A(n87), .B(addr[6]), .Y(n91) );
  NOR2X1 U55 ( .A(n7), .B(n1), .Y(n92) );
  CLKINVX1 U56 ( .A(n100), .Y(n8) );
  OA21XL U57 ( .A0(n1), .A1(n115), .B0(n120), .Y(n132) );
  AOI221XL U58 ( .A0(n13), .A1(n2), .B0(n15), .B1(addr[4]), .C0(n122), .Y(n126) );
  OAI22XL U59 ( .A0(n2), .A1(n14), .B0(addr[4]), .B1(n131), .Y(n122) );
  OAI211X1 U62 ( .A0(addr[2]), .A1(n99), .B0(n98), .C0(n97), .Y(dout[2]) );
  AOI221XL U63 ( .A0(addr[2]), .A1(n96), .B0(n1), .B1(n95), .C0(n94), .Y(n97)
         );
  AOI221XL U64 ( .A0(n91), .A1(n1), .B0(n90), .B1(n74), .C0(n89), .Y(n99) );
  OAI211X1 U65 ( .A0(n132), .A1(n131), .B0(n130), .C0(n129), .Y(dout[4]) );
  AOI222XL U66 ( .A0(n128), .A1(n4), .B0(n1), .B1(n127), .C0(n6), .C1(n15), 
        .Y(n129) );
  OAI211X1 U67 ( .A0(addr[1]), .A1(n114), .B0(n113), .C0(n112), .Y(dout[3]) );
  AOI221XL U68 ( .A0(n111), .A1(n9), .B0(n6), .B1(n13), .C0(n110), .Y(n112) );
  AOI2BB2XL U69 ( .B0(n102), .B1(n4), .A0N(n115), .A1N(n125), .Y(n113) );
  NAND4BX1 U70 ( .AN(n85), .B(n84), .C(n83), .D(n82), .Y(dout[1]) );
  AOI221XL U71 ( .A0(n12), .A1(n81), .B0(n3), .B1(n11), .C0(n80), .Y(n82) );
  AOI22X1 U72 ( .A0(n15), .A1(n77), .B0(n16), .B1(n76), .Y(n83) );
  CLKINVX3 U73 ( .A(addr[4]), .Y(n4) );
  CLKINVX3 U74 ( .A(addr[2]), .Y(n9) );
  CLKINVX3 U75 ( .A(n116), .Y(n10) );
  CLKINVX3 U76 ( .A(addr[1]), .Y(n14) );
  CLKINVX3 U77 ( .A(n105), .Y(n15) );
  CLKINVX3 U78 ( .A(n1), .Y(n74) );
  CLKINVX3 U79 ( .A(addr[6]), .Y(n75) );
endmodule


module crp_5 ( P, R, K_sub );
  output [1:32] P;
  input [1:32] R;
  input [1:48] K_sub;
  wire   n1;
  wire   [1:48] X;

  sbox1_5 u0 ( .addr(X[1:6]), .dout({P[9], P[17], P[23], P[31]}) );
  sbox2_5 u1 ( .addr({X[7], n1, X[9:12]}), .dout({P[13], P[28], P[2], P[18]})
         );
  sbox3_5 u2 ( .addr(X[13:18]), .dout({P[24], P[16], P[30], P[6]}) );
  sbox4_5 u3 ( .addr(X[19:24]), .dout({P[26], P[20], P[10], P[1]}) );
  sbox5_5 u4 ( .addr(X[25:30]), .dout({P[8], P[14], P[25], P[3]}) );
  sbox6_5 u5 ( .addr(X[31:36]), .dout({P[4], P[29], P[11], P[19]}) );
  sbox7_5 u6 ( .addr(X[37:42]), .dout({P[32], P[12], P[22], P[7]}) );
  sbox8_5 u7 ( .addr(X[43:48]), .dout({P[5], P[27], P[15], P[21]}) );
  XNOR2X1 U1 ( .A(R[5]), .B(K_sub[8]), .Y(X[8]) );
  INVX3 U2 ( .A(X[8]), .Y(n1) );
  XOR2X1 U3 ( .A(R[1]), .B(K_sub[2]), .Y(X[2]) );
  CLKXOR2X4 U4 ( .A(R[29]), .B(K_sub[42]), .Y(X[42]) );
  CLKXOR2X4 U5 ( .A(R[8]), .B(K_sub[11]), .Y(X[11]) );
  CLKXOR2X4 U6 ( .A(R[22]), .B(K_sub[33]), .Y(X[33]) );
  CLKXOR2X4 U7 ( .A(R[16]), .B(K_sub[25]), .Y(X[25]) );
  CLKXOR2X4 U8 ( .A(R[29]), .B(K_sub[44]), .Y(X[44]) );
  CLKXOR2X4 U9 ( .A(R[12]), .B(K_sub[19]), .Y(X[19]) );
  CLKXOR2X4 U10 ( .A(R[10]), .B(K_sub[15]), .Y(X[15]) );
  CLKXOR2X4 U11 ( .A(R[20]), .B(K_sub[31]), .Y(X[31]) );
  CLKXOR2X4 U12 ( .A(R[16]), .B(K_sub[23]), .Y(X[23]) );
  CLKXOR2X4 U13 ( .A(R[31]), .B(K_sub[46]), .Y(X[46]) );
  CLKXOR2X4 U14 ( .A(R[26]), .B(K_sub[39]), .Y(X[39]) );
  CLKXOR2X4 U15 ( .A(R[20]), .B(K_sub[29]), .Y(X[29]) );
  CLKXOR2X2 U16 ( .A(R[4]), .B(K_sub[5]), .Y(X[5]) );
  CLKXOR2X2 U17 ( .A(R[15]), .B(K_sub[22]), .Y(X[22]) );
  CLKXOR2X2 U18 ( .A(R[24]), .B(K_sub[35]), .Y(X[35]) );
  CLKXOR2X2 U19 ( .A(R[21]), .B(K_sub[30]), .Y(X[30]) );
  CLKXOR2X2 U20 ( .A(R[12]), .B(K_sub[17]), .Y(X[17]) );
  CLKXOR2X2 U21 ( .A(R[32]), .B(K_sub[1]), .Y(X[1]) );
  CLKXOR2X2 U22 ( .A(R[13]), .B(K_sub[20]), .Y(X[20]) );
  CLKXOR2X2 U23 ( .A(R[18]), .B(K_sub[27]), .Y(X[27]) );
  CLKXOR2X2 U24 ( .A(R[8]), .B(K_sub[13]), .Y(X[13]) );
  CLKXOR2X2 U25 ( .A(R[5]), .B(K_sub[6]), .Y(X[6]) );
  CLKXOR2X2 U26 ( .A(R[4]), .B(K_sub[7]), .Y(X[7]) );
  CLKXOR2X2 U27 ( .A(R[24]), .B(K_sub[37]), .Y(X[37]) );
  CLKXOR2X2 U28 ( .A(R[28]), .B(K_sub[43]), .Y(X[43]) );
  CLKXOR2X2 U29 ( .A(R[1]), .B(K_sub[48]), .Y(X[48]) );
  CLKXOR2X2 U30 ( .A(R[17]), .B(K_sub[24]), .Y(X[24]) );
  CLKXOR2X2 U31 ( .A(R[9]), .B(K_sub[12]), .Y(X[12]) );
  CLKXOR2X2 U32 ( .A(R[13]), .B(K_sub[18]), .Y(X[18]) );
  CLKXOR2X2 U33 ( .A(R[25]), .B(K_sub[36]), .Y(X[36]) );
  XOR2X1 U34 ( .A(R[23]), .B(K_sub[34]), .Y(X[34]) );
  XOR2X1 U35 ( .A(R[9]), .B(K_sub[14]), .Y(X[14]) );
  XOR2X1 U36 ( .A(R[30]), .B(K_sub[45]), .Y(X[45]) );
  XOR2X1 U37 ( .A(R[21]), .B(K_sub[32]), .Y(X[32]) );
  XOR2X1 U38 ( .A(R[25]), .B(K_sub[38]), .Y(X[38]) );
  XOR2X1 U39 ( .A(R[27]), .B(K_sub[40]), .Y(X[40]) );
  XOR2X1 U40 ( .A(R[3]), .B(K_sub[4]), .Y(X[4]) );
  XOR2X1 U41 ( .A(R[11]), .B(K_sub[16]), .Y(X[16]) );
  XOR2X1 U42 ( .A(R[7]), .B(K_sub[10]), .Y(X[10]) );
  XOR2X1 U43 ( .A(R[14]), .B(K_sub[21]), .Y(X[21]) );
  XOR2X1 U44 ( .A(R[6]), .B(K_sub[9]), .Y(X[9]) );
  XOR2X1 U45 ( .A(R[2]), .B(K_sub[3]), .Y(X[3]) );
  XOR2X1 U46 ( .A(R[28]), .B(K_sub[41]), .Y(X[41]) );
  XOR2X1 U47 ( .A(R[17]), .B(K_sub[26]), .Y(X[26]) );
  XOR2X1 U48 ( .A(R[32]), .B(K_sub[47]), .Y(X[47]) );
  XOR2X1 U49 ( .A(R[19]), .B(K_sub[28]), .Y(X[28]) );
endmodule


module sbox1_4 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127;

  OAI222X4 U13 ( .A0(addr[5]), .A1(n101), .B0(n1), .B1(n100), .C0(n99), .C1(n8), .Y(dout[3]) );
  OAI21X2 U42 ( .A0(n4), .A1(n112), .B0(n106), .Y(n123) );
  NAND2X2 U44 ( .A(addr[6]), .B(n13), .Y(n115) );
  NAND2X2 U48 ( .A(addr[1]), .B(n71), .Y(n114) );
  OAI22X2 U49 ( .A0(n72), .A1(n6), .B0(addr[5]), .B1(n120), .Y(n85) );
  NAND2X2 U50 ( .A(n3), .B(n72), .Y(n120) );
  NOR2X2 U51 ( .A(n72), .B(n3), .Y(n124) );
  NOR3X2 U55 ( .A(n2), .B(addr[6]), .C(n8), .Y(n102) );
  NOR2X2 U56 ( .A(n109), .B(n3), .Y(n93) );
  NAND2X2 U57 ( .A(addr[1]), .B(addr[6]), .Y(n109) );
  NAND2X2 U59 ( .A(n13), .B(n71), .Y(n112) );
  NOR2X1 U1 ( .A(n114), .B(n120), .Y(n104) );
  BUFX4 U2 ( .A(addr[4]), .Y(n2) );
  CLKBUFX3 U3 ( .A(addr[2]), .Y(n1) );
  OAI32X1 U4 ( .A0(n112), .A1(n2), .A2(n4), .B0(n115), .B1(n113), .Y(n80) );
  NOR2BXL U5 ( .AN(n118), .B(n1), .Y(n122) );
  CLKBUFX3 U6 ( .A(addr[2]), .Y(n4) );
  INVX3 U7 ( .A(addr[6]), .Y(n71) );
  OAI221X4 U8 ( .A0(n88), .A1(n6), .B0(addr[5]), .B1(n87), .C0(n86), .Y(
        dout[2]) );
  OAI221X4 U9 ( .A0(addr[5]), .A1(n127), .B0(n126), .B1(n6), .C0(n125), .Y(
        dout[4]) );
  OA21XL U10 ( .A0(n95), .A1(n115), .B0(n107), .Y(n119) );
  AOI222XL U11 ( .A0(n12), .A1(n1), .B0(n2), .B1(n110), .C0(n69), .C1(n8), .Y(
        n111) );
  AOI2BB2X1 U12 ( .B0(n2), .B1(n69), .A0N(addr[4]), .A1N(n115), .Y(n91) );
  BUFX4 U14 ( .A(addr[3]), .Y(n3) );
  CLKINVX1 U15 ( .A(n112), .Y(n12) );
  CLKINVX1 U16 ( .A(n113), .Y(n7) );
  NAND2BX1 U17 ( .AN(n104), .B(n119), .Y(n84) );
  CLKXOR2X2 U18 ( .A(n9), .B(n8), .Y(n90) );
  NOR2X1 U19 ( .A(n72), .B(n9), .Y(n118) );
  OAI21XL U20 ( .A0(n9), .A1(n114), .B0(n91), .Y(n92) );
  NAND2X1 U21 ( .A(n93), .B(n72), .Y(n107) );
  NAND2X1 U22 ( .A(n8), .B(n9), .Y(n113) );
  OAI211X1 U23 ( .A0(n72), .A1(n114), .B0(n108), .C0(n107), .Y(n89) );
  CLKINVX1 U24 ( .A(n109), .Y(n69) );
  NAND2X1 U25 ( .A(n124), .B(n11), .Y(n108) );
  CLKINVX1 U26 ( .A(n114), .Y(n70) );
  CLKINVX1 U27 ( .A(n115), .Y(n11) );
  CLKINVX1 U28 ( .A(n95), .Y(n5) );
  AO22X1 U29 ( .A0(n90), .A1(n11), .B0(n9), .B1(n123), .Y(n76) );
  OAI31X1 U30 ( .A0(n8), .A1(n3), .A2(n13), .B0(n103), .Y(n105) );
  AOI31XL U31 ( .A0(n13), .A1(n8), .A2(n2), .B0(n102), .Y(n103) );
  AOI211X1 U32 ( .A0(n10), .A1(n4), .B0(n117), .C0(n116), .Y(n126) );
  CLKINVX1 U33 ( .A(n108), .Y(n10) );
  AOI211X1 U34 ( .A0(n115), .A1(n114), .B0(n113), .C0(n2), .Y(n116) );
  OAI22X1 U35 ( .A0(n120), .A1(n112), .B0(n111), .B1(n9), .Y(n117) );
  AOI211X1 U36 ( .A0(n69), .A1(n118), .B0(n81), .C0(n80), .Y(n88) );
  OAI22X1 U37 ( .A0(n91), .A1(n8), .B0(n3), .B1(n106), .Y(n81) );
  CLKINVX3 U38 ( .A(addr[5]), .Y(n6) );
  NAND2X1 U39 ( .A(n3), .B(n6), .Y(n95) );
  NAND2X1 U40 ( .A(n70), .B(n1), .Y(n106) );
  XOR2X1 U41 ( .A(n82), .B(n2), .Y(n83) );
  NAND2X1 U43 ( .A(n1), .B(n3), .Y(n82) );
  OAI22XL U45 ( .A0(n3), .A1(n13), .B0(n9), .B1(n112), .Y(n94) );
  AOI211XL U46 ( .A0(n98), .A1(n9), .B0(n97), .C0(n104), .Y(n99) );
  OAI22XL U47 ( .A0(n96), .A1(n72), .B0(n95), .B1(n109), .Y(n97) );
  OAI22XL U52 ( .A0(n71), .A1(n6), .B0(n2), .B1(addr[1]), .Y(n98) );
  AOI221XL U53 ( .A0(n5), .A1(addr[6]), .B0(addr[5]), .B1(n94), .C0(n93), .Y(
        n96) );
  OAI21XL U54 ( .A0(addr[1]), .A1(n120), .B0(n119), .Y(n121) );
  AOI221XL U58 ( .A0(n12), .A1(n118), .B0(n93), .B1(n6), .C0(n75), .Y(n78) );
  OAI31X1 U60 ( .A0(n6), .A1(n2), .A2(n74), .B0(n73), .Y(n75) );
  OA21XL U61 ( .A0(n3), .A1(n71), .B0(n109), .Y(n74) );
  OAI21XL U62 ( .A0(n124), .A1(n85), .B0(n70), .Y(n73) );
  OAI21XL U63 ( .A0(n1), .A1(n13), .B0(n109), .Y(n110) );
  INVX4 U64 ( .A(n4), .Y(n8) );
  AOI222XL U65 ( .A0(n124), .A1(n123), .B0(n122), .B1(addr[6]), .C0(n1), .C1(
        n121), .Y(n125) );
  NOR4BBX1 U66 ( .AN(n107), .BN(n106), .C(n105), .D(n104), .Y(n127) );
  AOI222XL U67 ( .A0(n12), .A1(n90), .B0(n89), .B1(n8), .C0(n123), .C1(n72), 
        .Y(n101) );
  AOI2BB2XL U68 ( .B0(addr[5]), .B1(n92), .A0N(n120), .A1N(addr[1]), .Y(n100)
         );
  AOI32X1 U69 ( .A0(n4), .A1(n85), .A2(n12), .B0(n84), .B1(n8), .Y(n86) );
  AOI222XL U70 ( .A0(n124), .A1(n13), .B0(n83), .B1(addr[1]), .C0(n7), .C1(n71), .Y(n87) );
  OAI221X1 U71 ( .A0(n79), .A1(n6), .B0(n4), .B1(n78), .C0(n77), .Y(dout[1])
         );
  AOI32XL U72 ( .A0(addr[6]), .A1(n85), .A2(n1), .B0(n76), .B1(n6), .Y(n77) );
  AOI221X1 U73 ( .A0(n12), .A1(n90), .B0(n4), .B1(n93), .C0(n102), .Y(n79) );
  CLKINVX3 U74 ( .A(n3), .Y(n9) );
  CLKINVX3 U75 ( .A(addr[1]), .Y(n13) );
  CLKINVX3 U76 ( .A(n2), .Y(n72) );
endmodule


module sbox2_4 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147;

  NAND2X2 U55 ( .A(n2), .B(n16), .Y(n136) );
  NAND2X2 U57 ( .A(addr[2]), .B(n5), .Y(n104) );
  NAND2X2 U60 ( .A(addr[5]), .B(addr[2]), .Y(n132) );
  NOR2X2 U61 ( .A(n10), .B(n8), .Y(n101) );
  NAND2X2 U62 ( .A(n83), .B(n9), .Y(n146) );
  NAND2X2 U63 ( .A(n3), .B(n13), .Y(n124) );
  NAND2X2 U64 ( .A(addr[6]), .B(n83), .Y(n122) );
  NAND2X2 U67 ( .A(n3), .B(n2), .Y(n133) );
  AOI222XL U1 ( .A0(n15), .A1(n7), .B0(n88), .B1(n13), .C0(n140), .C1(n8), .Y(
        n89) );
  CLKINVX1 U2 ( .A(n121), .Y(n10) );
  CLKINVX1 U3 ( .A(addr[5]), .Y(n1) );
  INVX3 U4 ( .A(addr[5]), .Y(n5) );
  OAI211X4 U5 ( .A0(n147), .A1(n146), .B0(n145), .C0(n144), .Y(dout[4]) );
  NAND3XL U6 ( .A(n98), .B(n97), .C(n96), .Y(dout[1]) );
  NOR2X1 U7 ( .A(n104), .B(n2), .Y(n141) );
  NOR2X1 U8 ( .A(n124), .B(n2), .Y(n140) );
  CLKBUFX4 U9 ( .A(addr[4]), .Y(n2) );
  NAND2X1 U10 ( .A(addr[1]), .B(addr[6]), .Y(n121) );
  CLKINVX2 U11 ( .A(addr[1]), .Y(n83) );
  OAI221X1 U12 ( .A0(addr[1]), .A1(n136), .B0(n133), .B1(n83), .C0(n87), .Y(
        n95) );
  NAND2X4 U13 ( .A(addr[1]), .B(n9), .Y(n114) );
  INVX3 U14 ( .A(addr[6]), .Y(n9) );
  NAND2XL U15 ( .A(n102), .B(n16), .Y(n109) );
  AOI211XL U16 ( .A0(n6), .A1(n95), .B0(n94), .C0(n93), .Y(n96) );
  AOI2BB2X1 U17 ( .B0(n5), .B1(n12), .A0N(n104), .A1N(n136), .Y(n117) );
  NOR3BXL U18 ( .AN(n135), .B(n134), .C(n15), .Y(n147) );
  BUFX4 U19 ( .A(addr[3]), .Y(n3) );
  NAND2X1 U20 ( .A(n15), .B(n10), .Y(n113) );
  CLKINVX1 U21 ( .A(n146), .Y(n8) );
  CLKINVX1 U22 ( .A(n115), .Y(n15) );
  CLKINVX1 U23 ( .A(n122), .Y(n11) );
  OAI31X1 U24 ( .A0(n124), .A1(n9), .A2(n5), .B0(n123), .Y(n128) );
  OAI21XL U25 ( .A0(n5), .A1(n83), .B0(n140), .Y(n123) );
  OAI22X1 U26 ( .A0(n122), .A1(n124), .B0(n101), .B1(n132), .Y(n84) );
  INVX1 U27 ( .A(n114), .Y(n7) );
  OAI22X1 U28 ( .A0(n122), .A1(n16), .B0(n82), .B1(n121), .Y(n129) );
  NAND3X1 U29 ( .A(n82), .B(n5), .C(n83), .Y(n111) );
  NAND2X1 U30 ( .A(n16), .B(n82), .Y(n115) );
  OAI21XL U31 ( .A0(n13), .A1(n133), .B0(n135), .Y(n85) );
  OAI22XL U32 ( .A0(n117), .A1(n146), .B0(n116), .B1(n132), .Y(n118) );
  AOI222XL U33 ( .A0(n7), .A1(n115), .B0(n81), .B1(n9), .C0(n15), .C1(n8), .Y(
        n116) );
  CLKINVX1 U34 ( .A(n104), .Y(n4) );
  OAI2BB2XL U35 ( .B0(n114), .B1(n135), .A0N(n126), .A1N(n81), .Y(n106) );
  OAI21XL U36 ( .A0(n112), .A1(n114), .B0(n111), .Y(n120) );
  OAI21XL U37 ( .A0(n133), .A1(n114), .B0(n113), .Y(n119) );
  CLKINVX1 U38 ( .A(n124), .Y(n12) );
  CLKINVX1 U39 ( .A(n136), .Y(n14) );
  CLKINVX1 U40 ( .A(n133), .Y(n81) );
  CLKINVX1 U41 ( .A(n132), .Y(n6) );
  AOI2BB1X1 U42 ( .A0N(n126), .A1N(n125), .B0(n136), .Y(n127) );
  OAI22XL U43 ( .A0(n104), .A1(n114), .B0(n101), .B1(n132), .Y(n102) );
  AO21XL U44 ( .A0(n13), .A1(n14), .B0(n141), .Y(n86) );
  AO21X1 U45 ( .A0(n16), .A1(n4), .B0(n140), .Y(n142) );
  NAND3X1 U46 ( .A(n13), .B(n82), .C(addr[5]), .Y(n135) );
  OAI22X1 U47 ( .A0(addr[5]), .A1(n121), .B0(n122), .B1(n5), .Y(n126) );
  AOI2BB1X1 U48 ( .A0N(n3), .A1N(n1), .B0(n14), .Y(n112) );
  NOR3X1 U49 ( .A(addr[1]), .B(addr[2]), .C(n5), .Y(n125) );
  AOI2BB1XL U50 ( .A0N(n92), .A1N(n91), .B0(addr[5]), .Y(n93) );
  OAI22XL U51 ( .A0(n117), .A1(n114), .B0(n89), .B1(n1), .Y(n94) );
  OAI31XL U52 ( .A0(n114), .A1(n2), .A2(n16), .B0(n90), .Y(n91) );
  OAI21XL U53 ( .A0(n81), .A1(n12), .B0(n11), .Y(n90) );
  NAND2X1 U54 ( .A(n7), .B(n2), .Y(n137) );
  OAI31XL U56 ( .A0(n101), .A1(n3), .A2(addr[2]), .B0(n113), .Y(n92) );
  OAI211X1 U58 ( .A0(n139), .A1(n5), .B0(n138), .C0(n137), .Y(n143) );
  NAND3X1 U59 ( .A(n82), .B(n5), .C(addr[6]), .Y(n138) );
  AOI2BB2X1 U65 ( .B0(n11), .B1(n16), .A0N(n83), .A1N(n136), .Y(n139) );
  OAI22XL U66 ( .A0(addr[5]), .A1(n133), .B0(n3), .B1(n132), .Y(n134) );
  OAI2BB2XL U68 ( .B0(n112), .B1(n122), .A0N(n1), .A1N(n99), .Y(n100) );
  OAI211X1 U69 ( .A0(n146), .A1(n2), .B0(n137), .C0(n113), .Y(n99) );
  NAND3X1 U70 ( .A(n11), .B(n82), .C(n3), .Y(n87) );
  AOI2BB2XL U71 ( .B0(n3), .B1(n105), .A0N(n137), .A1N(n132), .Y(n108) );
  OAI211XL U72 ( .A0(n104), .A1(n146), .B0(n103), .C0(n111), .Y(n105) );
  NAND3XL U73 ( .A(addr[5]), .B(n82), .C(n10), .Y(n103) );
  OAI22XL U74 ( .A0(n3), .A1(n114), .B0(n9), .B1(n115), .Y(n88) );
  NAND4X1 U75 ( .A(n110), .B(n109), .C(n108), .D(n107), .Y(dout[2]) );
  AOI32XL U76 ( .A0(addr[1]), .A1(addr[2]), .A2(n14), .B0(n100), .B1(n13), .Y(
        n110) );
  AOI221XL U77 ( .A0(n125), .A1(addr[4]), .B0(n141), .B1(n11), .C0(n106), .Y(
        n107) );
  AOI33XL U78 ( .A0(n11), .A1(n4), .A2(n2), .B0(n6), .B1(n146), .B2(n3), .Y(
        n145) );
  AOI222XL U79 ( .A0(n143), .A1(n13), .B0(n10), .B1(n142), .C0(n7), .C1(n141), 
        .Y(n144) );
  AOI32XL U80 ( .A0(n4), .A1(n83), .A2(n15), .B0(n8), .B1(n86), .Y(n97) );
  AOI22X1 U81 ( .A0(n10), .A1(n85), .B0(n2), .B1(n84), .Y(n98) );
  NAND2X1 U82 ( .A(n131), .B(n130), .Y(dout[3]) );
  AOI221XL U83 ( .A0(n120), .A1(n13), .B0(addr[2]), .B1(n119), .C0(n118), .Y(
        n131) );
  AOI211X1 U84 ( .A0(n4), .A1(n129), .B0(n128), .C0(n127), .Y(n130) );
  CLKINVX3 U85 ( .A(addr[2]), .Y(n13) );
  CLKINVX3 U86 ( .A(n3), .Y(n16) );
  CLKINVX3 U87 ( .A(n2), .Y(n82) );
endmodule


module sbox3_4 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134;

  NOR2X2 U35 ( .A(n78), .B(addr[3]), .Y(n109) );
  NOR2X2 U50 ( .A(addr[1]), .B(addr[6]), .Y(n108) );
  NOR2X2 U52 ( .A(n11), .B(n3), .Y(n88) );
  NOR2X2 U56 ( .A(n11), .B(n12), .Y(n95) );
  NOR2X1 U1 ( .A(n78), .B(n11), .Y(n107) );
  OAI221X1 U2 ( .A0(n125), .A1(n78), .B0(n4), .B1(addr[1]), .C0(n76), .Y(n105)
         );
  INVXL U3 ( .A(n2), .Y(n1) );
  NOR2X1 U4 ( .A(n17), .B(n4), .Y(n92) );
  NOR2X1 U5 ( .A(n8), .B(n4), .Y(n122) );
  NOR2X1 U6 ( .A(n76), .B(n4), .Y(n96) );
  CLKBUFX3 U7 ( .A(addr[2]), .Y(n4) );
  INVX1 U8 ( .A(addr[2]), .Y(n2) );
  NOR2X1 U9 ( .A(n4), .B(n3), .Y(n111) );
  BUFX4 U10 ( .A(addr[4]), .Y(n3) );
  OAI33X1 U11 ( .A0(n8), .A1(n126), .A2(n12), .B0(n78), .B1(n95), .B2(n120), 
        .Y(n80) );
  INVX3 U12 ( .A(n4), .Y(n12) );
  OAI221X1 U13 ( .A0(addr[5]), .A1(n91), .B0(n90), .B1(n77), .C0(n89), .Y(
        dout[1]) );
  NOR2X4 U14 ( .A(n18), .B(n79), .Y(n125) );
  NOR2X4 U15 ( .A(addr[3]), .B(n3), .Y(n131) );
  NOR2X4 U16 ( .A(n79), .B(addr[6]), .Y(n126) );
  INVX3 U17 ( .A(addr[1]), .Y(n79) );
  NAND2XL U18 ( .A(n95), .B(n125), .Y(n133) );
  OAI211XL U19 ( .A0(n3), .A1(n13), .B0(n129), .C0(n128), .Y(n130) );
  NAND4XL U20 ( .A(n115), .B(n114), .C(n113), .D(n112), .Y(n116) );
  CLKINVX1 U21 ( .A(n133), .Y(n10) );
  INVX1 U22 ( .A(n125), .Y(n15) );
  CLKINVX1 U23 ( .A(n107), .Y(n6) );
  NAND2X1 U24 ( .A(n17), .B(n19), .Y(n123) );
  CLKINVX1 U25 ( .A(n87), .Y(n19) );
  CLKINVX1 U26 ( .A(n121), .Y(n5) );
  CLKINVX1 U27 ( .A(n120), .Y(n16) );
  CLKINVX1 U28 ( .A(n115), .Y(n9) );
  CLKINVX1 U29 ( .A(n108), .Y(n76) );
  NOR2X1 U30 ( .A(n17), .B(n12), .Y(n104) );
  NOR2X1 U31 ( .A(n15), .B(n12), .Y(n110) );
  INVX1 U32 ( .A(n126), .Y(n20) );
  AOI21X1 U33 ( .A0(n11), .A1(n12), .B0(n95), .Y(n121) );
  OAI21XL U34 ( .A0(n111), .A1(n131), .B0(n125), .Y(n83) );
  CLKINVX1 U36 ( .A(n82), .Y(n17) );
  NOR2X1 U37 ( .A(n20), .B(n78), .Y(n87) );
  NOR2X1 U38 ( .A(n125), .B(n108), .Y(n120) );
  OAI21XL U39 ( .A0(n110), .A1(n92), .B0(n131), .Y(n101) );
  NAND2X1 U40 ( .A(n104), .B(n88), .Y(n115) );
  CLKINVX1 U41 ( .A(n88), .Y(n8) );
  CLKINVX1 U42 ( .A(n92), .Y(n13) );
  CLKINVX1 U43 ( .A(n111), .Y(n14) );
  CLKINVX1 U44 ( .A(n122), .Y(n7) );
  OR2X1 U45 ( .A(n104), .B(n96), .Y(n127) );
  OAI221X1 U46 ( .A0(n20), .A1(n14), .B0(n12), .B1(n19), .C0(n94), .Y(n99) );
  AOI221XL U47 ( .A0(n96), .A1(n3), .B0(n93), .B1(n78), .C0(n10), .Y(n94) );
  OAI21XL U48 ( .A0(n12), .A1(n76), .B0(n13), .Y(n93) );
  XNOR2X1 U49 ( .A(addr[5]), .B(addr[3]), .Y(n103) );
  CLKINVX1 U51 ( .A(addr[5]), .Y(n77) );
  OAI221X1 U53 ( .A0(n76), .A1(n14), .B0(n15), .B1(n8), .C0(n106), .Y(n117) );
  AOI221XL U54 ( .A0(addr[3]), .A1(n105), .B0(n104), .B1(n131), .C0(n10), .Y(
        n106) );
  CLKINVX1 U55 ( .A(addr[6]), .Y(n18) );
  NAND3X1 U57 ( .A(n4), .B(n79), .C(n109), .Y(n114) );
  NOR2X1 U58 ( .A(n18), .B(addr[1]), .Y(n82) );
  AOI32XL U59 ( .A0(n12), .A1(n11), .A2(n125), .B0(n124), .B1(n18), .Y(n129)
         );
  AOI22XL U60 ( .A0(n3), .A1(n127), .B0(n126), .B1(n131), .Y(n128) );
  OAI22XL U61 ( .A0(n3), .A1(n2), .B0(n4), .B1(n6), .Y(n124) );
  AOI222XL U62 ( .A0(n111), .A1(n126), .B0(n110), .B1(n11), .C0(n109), .C1(
        n108), .Y(n112) );
  OAI211XL U63 ( .A0(n107), .A1(n131), .B0(n2), .C0(addr[6]), .Y(n113) );
  OAI21XL U64 ( .A0(n1), .A1(addr[1]), .B0(n20), .Y(n81) );
  AOI221XL U65 ( .A0(n87), .A1(n11), .B0(n88), .B1(n126), .C0(n86), .Y(n90) );
  OAI211X1 U66 ( .A0(n85), .A1(n12), .B0(n84), .C0(n83), .Y(n86) );
  AOI222XL U67 ( .A0(n82), .A1(n11), .B0(n108), .B1(n107), .C0(n131), .C1(n79), 
        .Y(n85) );
  OAI21XL U68 ( .A0(n92), .A1(n10), .B0(addr[4]), .Y(n84) );
  AOI221XL U69 ( .A0(n126), .A1(n5), .B0(addr[3]), .B1(n127), .C0(n97), .Y(n98) );
  OAI22X1 U70 ( .A0(n15), .A1(n7), .B0(n6), .B1(n17), .Y(n97) );
  OAI211X1 U71 ( .A0(n76), .A1(n7), .B0(n119), .C0(n118), .Y(dout[3]) );
  AOI32XL U72 ( .A0(n126), .A1(n4), .A2(n103), .B0(n109), .B1(n110), .Y(n119)
         );
  AOI22XL U73 ( .A0(n117), .A1(n77), .B0(addr[5]), .B1(n116), .Y(n118) );
  AOI221XL U74 ( .A0(n122), .A1(n126), .B0(n96), .B1(n109), .C0(n9), .Y(n89)
         );
  AOI221XL U75 ( .A0(n131), .A1(n81), .B0(n95), .B1(n123), .C0(n80), .Y(n91)
         );
  NAND4X1 U76 ( .A(n102), .B(n114), .C(n101), .D(n100), .Y(dout[2]) );
  NAND3XL U77 ( .A(n3), .B(n125), .C(n103), .Y(n102) );
  AOI2BB2XL U78 ( .B0(addr[5]), .B1(n99), .A0N(addr[5]), .A1N(n98), .Y(n100)
         );
  OAI221X1 U79 ( .A0(n134), .A1(n77), .B0(n3), .B1(n133), .C0(n132), .Y(
        dout[4]) );
  AOI32XL U80 ( .A0(n131), .A1(n18), .A2(n1), .B0(n130), .B1(n77), .Y(n132) );
  AOI222XL U81 ( .A0(n5), .A1(n123), .B0(n122), .B1(addr[1]), .C0(n121), .C1(
        n16), .Y(n134) );
  CLKINVX3 U82 ( .A(addr[3]), .Y(n11) );
  CLKINVX3 U83 ( .A(n3), .Y(n78) );
endmodule


module sbox4_4 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126;

  OAI32X4 U12 ( .A0(n6), .A1(n2), .A2(addr[2]), .B0(n5), .B1(n108), .Y(n123)
         );
  OAI222X4 U20 ( .A0(addr[2]), .A1(n92), .B0(n106), .B1(n91), .C0(n90), .C1(
        n72), .Y(dout[2]) );
  OAI222X4 U33 ( .A0(addr[4]), .A1(n106), .B0(n16), .B1(n108), .C0(n2), .C1(
        n118), .Y(n83) );
  NAND2X2 U34 ( .A(addr[4]), .B(n2), .Y(n108) );
  NOR2X2 U43 ( .A(n71), .B(addr[4]), .Y(n113) );
  NOR2X2 U45 ( .A(n5), .B(n2), .Y(n111) );
  NAND2X2 U51 ( .A(n16), .B(n11), .Y(n118) );
  NOR2X2 U52 ( .A(n15), .B(addr[5]), .Y(n97) );
  NAND2X2 U53 ( .A(addr[6]), .B(addr[1]), .Y(n85) );
  NAND2X2 U54 ( .A(addr[1]), .B(n11), .Y(n116) );
  NOR2X2 U55 ( .A(n115), .B(n5), .Y(n121) );
  NAND2X2 U56 ( .A(n71), .B(n15), .Y(n115) );
  NAND2X2 U57 ( .A(addr[5]), .B(n15), .Y(n96) );
  NAND2X2 U58 ( .A(addr[6]), .B(n16), .Y(n106) );
  OAI222X1 U1 ( .A0(n6), .A1(n85), .B0(n97), .B1(n116), .C0(n15), .C1(n118), 
        .Y(n73) );
  CLKINVX1 U2 ( .A(n116), .Y(n10) );
  CLKINVX1 U3 ( .A(n71), .Y(n1) );
  CLKBUFX3 U4 ( .A(addr[3]), .Y(n2) );
  OAI31X4 U5 ( .A0(n118), .A1(n5), .A2(n15), .B0(n117), .Y(n119) );
  OAI221X1 U6 ( .A0(addr[2]), .A1(n80), .B0(n118), .B1(n105), .C0(n79), .Y(
        dout[1]) );
  INVX4 U7 ( .A(addr[5]), .Y(n5) );
  OAI31X1 U8 ( .A0(n108), .A1(addr[5]), .A2(n12), .B0(n107), .Y(n109) );
  AOI222XL U9 ( .A0(n15), .A1(n11), .B0(n113), .B1(n16), .C0(addr[1]), .C1(n71), .Y(n114) );
  OAI222X1 U10 ( .A0(addr[1]), .A1(n84), .B0(n85), .B1(n74), .C0(n71), .C1(
        n107), .Y(n75) );
  NAND2XL U11 ( .A(n1), .B(addr[5]), .Y(n84) );
  AOI211XL U13 ( .A0(n83), .A1(n5), .B0(n82), .C0(n4), .Y(n92) );
  NAND2XL U14 ( .A(n15), .B(n5), .Y(n74) );
  CLKINVX1 U15 ( .A(n118), .Y(n8) );
  CLKINVX1 U16 ( .A(n115), .Y(n14) );
  CLKINVX1 U17 ( .A(n112), .Y(n9) );
  OAI21X1 U18 ( .A0(n10), .A1(n12), .B0(n72), .Y(n112) );
  AOI22X1 U19 ( .A0(n13), .A1(n111), .B0(n12), .B1(n113), .Y(n93) );
  OAI211X1 U21 ( .A0(n16), .A1(n115), .B0(n93), .C0(n3), .Y(n94) );
  CLKINVX1 U22 ( .A(n85), .Y(n13) );
  NAND2X1 U23 ( .A(n97), .B(n71), .Y(n105) );
  NAND2X1 U24 ( .A(n113), .B(n8), .Y(n98) );
  NAND2X1 U25 ( .A(n10), .B(n97), .Y(n107) );
  NAND2X1 U26 ( .A(n118), .B(n85), .Y(n110) );
  OAI21XL U27 ( .A0(n14), .A1(n5), .B0(n108), .Y(n95) );
  CLKINVX1 U28 ( .A(n84), .Y(n7) );
  CLKINVX1 U29 ( .A(addr[2]), .Y(n72) );
  OAI31X1 U30 ( .A0(n15), .A1(addr[6]), .A2(n5), .B0(n87), .Y(n88) );
  OAI21XL U31 ( .A0(n113), .A1(n6), .B0(n13), .Y(n87) );
  OAI211X1 U32 ( .A0(n76), .A1(n15), .B0(n98), .C0(n3), .Y(n77) );
  AOI222XL U35 ( .A0(addr[5]), .A1(addr[6]), .B0(n111), .B1(addr[1]), .C0(n12), 
        .C1(n2), .Y(n76) );
  NAND3XL U36 ( .A(n13), .B(n71), .C(addr[4]), .Y(n117) );
  OAI22XL U37 ( .A0(n116), .A1(n115), .B0(n1), .B1(n112), .Y(n78) );
  CLKINVX3 U38 ( .A(addr[4]), .Y(n15) );
  OAI2BB2XL U39 ( .B0(n115), .B1(n106), .A0N(n5), .A1N(n86), .Y(n89) );
  OAI221XL U40 ( .A0(n116), .A1(addr[4]), .B0(n108), .B1(addr[1]), .C0(n117), 
        .Y(n86) );
  CLKINVX1 U41 ( .A(addr[6]), .Y(n11) );
  CLKINVX1 U42 ( .A(n81), .Y(n4) );
  OAI21XL U44 ( .A0(n96), .A1(n118), .B0(n93), .Y(n82) );
  NAND3X1 U46 ( .A(n101), .B(n100), .C(n99), .Y(n102) );
  AOI32X1 U47 ( .A0(n96), .A1(n71), .A2(n10), .B0(n13), .B1(n95), .Y(n101) );
  AOI2BB2XL U48 ( .B0(n16), .B1(n121), .A0N(n98), .A1N(addr[5]), .Y(n99) );
  OAI21XL U49 ( .A0(n97), .A1(n6), .B0(n12), .Y(n100) );
  AOI2BB2XL U50 ( .B0(n12), .B1(n123), .A0N(n122), .A1N(n72), .Y(n124) );
  AOI211XL U59 ( .A0(n12), .A1(n121), .B0(n120), .C0(n119), .Y(n122) );
  OAI22XL U60 ( .A0(n116), .A1(n115), .B0(addr[5]), .B1(n114), .Y(n120) );
  CLKINVX1 U61 ( .A(n75), .Y(n3) );
  AOI32XL U62 ( .A0(n10), .A1(n96), .A2(n1), .B0(addr[1]), .B1(n121), .Y(n81)
         );
  AOI222XL U63 ( .A0(n12), .A1(n6), .B0(n121), .B1(n116), .C0(n2), .C1(n73), 
        .Y(n80) );
  AOI22XL U64 ( .A0(n78), .A1(n5), .B0(addr[2]), .B1(n77), .Y(n79) );
  NAND2XL U65 ( .A(n111), .B(addr[4]), .Y(n91) );
  AOI211X1 U66 ( .A0(n7), .A1(n110), .B0(n89), .C0(n88), .Y(n90) );
  OAI211X1 U67 ( .A0(n106), .A1(n105), .B0(n104), .C0(n103), .Y(dout[3]) );
  AOI32X1 U68 ( .A0(n2), .A1(n6), .A2(n10), .B0(n94), .B1(n72), .Y(n104) );
  AOI22XL U69 ( .A0(addr[2]), .A1(n102), .B0(n8), .B1(n123), .Y(n103) );
  OAI211X1 U70 ( .A0(addr[2]), .A1(n126), .B0(n125), .C0(n124), .Y(dout[4]) );
  AOI32X1 U71 ( .A0(n13), .A1(n6), .A2(n2), .B0(n9), .B1(n7), .Y(n125) );
  AOI221XL U72 ( .A0(n8), .A1(n111), .B0(n14), .B1(n110), .C0(n109), .Y(n126)
         );
  CLKINVX3 U73 ( .A(n96), .Y(n6) );
  CLKINVX3 U74 ( .A(n106), .Y(n12) );
  CLKINVX3 U75 ( .A(addr[1]), .Y(n16) );
  CLKINVX3 U76 ( .A(n2), .Y(n71) );
endmodule


module sbox5_4 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121;

  OAI222X4 U18 ( .A0(addr[3]), .A1(n106), .B0(n68), .B1(n90), .C0(n70), .C1(n8), .Y(n93) );
  OAI22X2 U40 ( .A0(addr[5]), .A1(n106), .B0(n69), .B1(n114), .Y(n116) );
  NOR2X2 U41 ( .A(n3), .B(addr[3]), .Y(n102) );
  NAND2X2 U45 ( .A(addr[6]), .B(n8), .Y(n114) );
  NAND2X2 U50 ( .A(n8), .B(n68), .Y(n110) );
  NAND2X2 U52 ( .A(addr[1]), .B(n68), .Y(n113) );
  NAND2X2 U54 ( .A(addr[1]), .B(addr[6]), .Y(n106) );
  NAND2X2 U55 ( .A(addr[3]), .B(n70), .Y(n121) );
  CLKINVX1 U1 ( .A(addr[5]), .Y(n1) );
  AOI221XL U2 ( .A0(n93), .A1(n1), .B0(n9), .B1(n13), .C0(n92), .Y(n105) );
  INVX3 U3 ( .A(addr[5]), .Y(n69) );
  OAI221X4 U4 ( .A0(n111), .A1(n110), .B0(n121), .B1(n114), .C0(n109), .Y(n112) );
  OAI221X4 U5 ( .A0(n70), .A1(n114), .B0(n69), .B1(n113), .C0(n120), .Y(n115)
         );
  OAI221X4 U6 ( .A0(n107), .A1(n121), .B0(n111), .B1(n113), .C0(n85), .Y(n86)
         );
  OAI31X1 U7 ( .A0(n14), .A1(addr[5]), .A2(addr[1]), .B0(n81), .Y(n73) );
  OAI32X1 U8 ( .A0(n114), .A1(addr[5]), .A2(n3), .B0(n15), .B1(n107), .Y(n79)
         );
  AOI32XL U9 ( .A0(n13), .A1(n98), .A2(n11), .B0(n2), .B1(n73), .Y(n77) );
  CLKBUFX3 U10 ( .A(addr[4]), .Y(n2) );
  CLKINVX1 U11 ( .A(n81), .Y(n4) );
  NAND2X1 U12 ( .A(n5), .B(n13), .Y(n81) );
  CLKINVX1 U13 ( .A(n110), .Y(n7) );
  CLKXOR2X2 U14 ( .A(n14), .B(n69), .Y(n94) );
  AOI2BB1X1 U15 ( .A0N(n70), .A1N(n1), .B0(n13), .Y(n111) );
  NOR2X1 U16 ( .A(n121), .B(n69), .Y(n91) );
  NOR2BX1 U17 ( .AN(n116), .B(n90), .Y(n83) );
  NAND2X1 U19 ( .A(n7), .B(n69), .Y(n120) );
  CLKINVX1 U20 ( .A(n113), .Y(n11) );
  NAND2X1 U21 ( .A(n11), .B(n69), .Y(n107) );
  CLKINVX1 U22 ( .A(n121), .Y(n15) );
  OAI31X1 U23 ( .A0(n12), .A1(n13), .A2(n113), .B0(n99), .Y(n72) );
  CLKINVX1 U24 ( .A(n106), .Y(n9) );
  OAI2BB2XL U25 ( .B0(n1), .B1(n113), .A0N(n98), .A1N(n5), .Y(n101) );
  CLKINVX1 U26 ( .A(n114), .Y(n5) );
  CLKINVX1 U27 ( .A(n90), .Y(n16) );
  CLKINVX1 U28 ( .A(addr[1]), .Y(n8) );
  CLKINVX1 U29 ( .A(addr[3]), .Y(n14) );
  CLKINVX1 U30 ( .A(addr[6]), .Y(n68) );
  AOI211X1 U31 ( .A0(n91), .A1(addr[1]), .B0(n80), .C0(n79), .Y(n89) );
  OAI2BB2XL U32 ( .B0(n111), .B1(n106), .A0N(n94), .A1N(n7), .Y(n80) );
  AOI211X1 U33 ( .A0(n102), .A1(n84), .B0(n83), .C0(n82), .Y(n85) );
  OAI21XL U34 ( .A0(n68), .A1(n1), .B0(n106), .Y(n84) );
  NOR3XL U35 ( .A(n94), .B(n3), .C(n110), .Y(n82) );
  AOI222XL U36 ( .A0(n9), .A1(n16), .B0(addr[5]), .B1(n108), .C0(n10), .C1(n70), .Y(n109) );
  CLKINVX1 U37 ( .A(n107), .Y(n10) );
  OAI21XL U38 ( .A0(addr[6]), .A1(addr[3]), .B0(n106), .Y(n108) );
  NAND2X1 U39 ( .A(addr[3]), .B(n3), .Y(n90) );
  NAND2X1 U42 ( .A(n2), .B(addr[5]), .Y(n98) );
  NAND2X1 U43 ( .A(n3), .B(n14), .Y(n97) );
  OAI21XL U44 ( .A0(addr[1]), .A1(n97), .B0(n96), .Y(n103) );
  AOI33XL U46 ( .A0(n3), .A1(n95), .A2(addr[5]), .B0(n94), .B1(n70), .B2(
        addr[1]), .Y(n96) );
  OAI21XL U47 ( .A0(n8), .A1(n14), .B0(n114), .Y(n95) );
  OAI21XL U48 ( .A0(addr[6]), .A1(n121), .B0(n99), .Y(n100) );
  NAND2X1 U49 ( .A(n71), .B(n7), .Y(n99) );
  XOR2X1 U51 ( .A(n12), .B(n3), .Y(n71) );
  AOI2BB2XL U53 ( .B0(n102), .B1(n116), .A0N(n2), .A1N(n75), .Y(n76) );
  AOI211X1 U56 ( .A0(n6), .A1(n3), .B0(n74), .C0(n83), .Y(n75) );
  AO22XL U57 ( .A0(n11), .A1(n15), .B0(addr[6]), .B1(n102), .Y(n74) );
  CLKINVX1 U58 ( .A(n120), .Y(n6) );
  CLKINVX1 U59 ( .A(n2), .Y(n12) );
  AO22XL U60 ( .A0(n11), .A1(n16), .B0(addr[6]), .B1(n91), .Y(n92) );
  AOI222XL U61 ( .A0(n116), .A1(n70), .B0(addr[3]), .B1(n115), .C0(n11), .C1(
        n13), .Y(n117) );
  OAI221X1 U62 ( .A0(n2), .A1(n105), .B0(n110), .B1(n121), .C0(n104), .Y(
        dout[3]) );
  AOI222XL U63 ( .A0(n2), .A1(n103), .B0(n102), .B1(n101), .C0(n100), .C1(n1), 
        .Y(n104) );
  OAI211X1 U64 ( .A0(n2), .A1(n89), .B0(n88), .C0(n87), .Y(dout[2]) );
  AOI33XL U65 ( .A0(n15), .A1(n98), .A2(n5), .B0(n3), .B1(n94), .B2(n7), .Y(
        n88) );
  AOI222XL U66 ( .A0(n4), .A1(n69), .B0(n2), .B1(n86), .C0(n91), .C1(n9), .Y(
        n87) );
  OAI211X1 U67 ( .A0(n78), .A1(n69), .B0(n77), .C0(n76), .Y(dout[1]) );
  AOI221XL U68 ( .A0(n15), .A1(addr[1]), .B0(n9), .B1(n13), .C0(n72), .Y(n78)
         );
  OAI211X1 U69 ( .A0(n121), .A1(n120), .B0(n119), .C0(n118), .Y(dout[4]) );
  AOI32XL U70 ( .A0(n13), .A1(n114), .A2(addr[5]), .B0(n2), .B1(n112), .Y(n119) );
  AOI2BB2X1 U71 ( .B0(n4), .B1(n69), .A0N(n2), .A1N(n117), .Y(n118) );
  BUFX4 U72 ( .A(addr[2]), .Y(n3) );
  CLKINVX3 U73 ( .A(n97), .Y(n13) );
  CLKINVX3 U74 ( .A(n3), .Y(n70) );
endmodule


module sbox6_4 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147;

  NAND2X2 U39 ( .A(n138), .B(addr[3]), .Y(n147) );
  NOR2X2 U47 ( .A(n84), .B(n12), .Y(n138) );
  NOR2X2 U50 ( .A(n85), .B(n4), .Y(n119) );
  NOR2X2 U58 ( .A(n81), .B(n85), .Y(n125) );
  NAND2X2 U61 ( .A(n97), .B(n103), .Y(n112) );
  NOR2X2 U62 ( .A(n83), .B(addr[1]), .Y(n103) );
  NOR2X2 U63 ( .A(n81), .B(addr[3]), .Y(n97) );
  NAND2X2 U64 ( .A(n117), .B(n131), .Y(n140) );
  NOR2X2 U65 ( .A(n5), .B(addr[3]), .Y(n131) );
  NOR2X2 U66 ( .A(n13), .B(addr[6]), .Y(n117) );
  NOR2X1 U1 ( .A(n84), .B(addr[3]), .Y(n102) );
  CLKINVX1 U2 ( .A(addr[3]), .Y(n1) );
  INVX3 U3 ( .A(addr[3]), .Y(n85) );
  CLKINVX1 U4 ( .A(n81), .Y(n2) );
  INVX4 U5 ( .A(n4), .Y(n81) );
  CLKBUFX3 U6 ( .A(addr[4]), .Y(n4) );
  CLKINVX1 U7 ( .A(n84), .Y(n3) );
  OAI222X1 U8 ( .A0(n91), .A1(n7), .B0(n5), .B1(n18), .C0(addr[5]), .C1(n82), 
        .Y(n92) );
  BUFX4 U9 ( .A(addr[2]), .Y(n5) );
  OAI221X1 U10 ( .A0(n83), .A1(n17), .B0(n85), .B1(n10), .C0(n86), .Y(n90) );
  INVX3 U11 ( .A(n96), .Y(n10) );
  NOR2X4 U12 ( .A(addr[1]), .B(addr[6]), .Y(n130) );
  OAI221X4 U13 ( .A0(n123), .A1(n15), .B0(n12), .B1(n7), .C0(n9), .Y(n124) );
  NOR2X4 U14 ( .A(n5), .B(addr[5]), .Y(n143) );
  INVX1 U15 ( .A(n130), .Y(n16) );
  CLKINVX1 U16 ( .A(n125), .Y(n17) );
  NAND2X1 U17 ( .A(n16), .B(n10), .Y(n105) );
  INVXL U18 ( .A(n121), .Y(n6) );
  CLKINVX1 U19 ( .A(n138), .Y(n11) );
  AOI211X1 U20 ( .A0(n7), .A1(n85), .B0(n131), .C0(n143), .Y(n121) );
  CLKINVX1 U21 ( .A(n117), .Y(n12) );
  CLKINVX1 U22 ( .A(n119), .Y(n82) );
  NOR2X1 U23 ( .A(n10), .B(n123), .Y(n144) );
  NOR2X1 U24 ( .A(n13), .B(n83), .Y(n96) );
  CLKINVX1 U25 ( .A(n103), .Y(n15) );
  OAI211X1 U26 ( .A0(n16), .A1(n17), .B0(n104), .C0(n112), .Y(n108) );
  OAI21XL U27 ( .A0(n103), .A1(n117), .B0(n102), .Y(n104) );
  OAI21XL U28 ( .A0(n132), .A1(n83), .B0(n1), .Y(n86) );
  AOI21X1 U29 ( .A0(n81), .A1(n102), .B0(n125), .Y(n91) );
  OAI2BB2XL U30 ( .B0(n143), .B1(n16), .A0N(n143), .A1N(n117), .Y(n118) );
  CLKINVX1 U31 ( .A(n122), .Y(n9) );
  CLKINVX1 U32 ( .A(n126), .Y(n14) );
  CLKINVX1 U33 ( .A(n97), .Y(n18) );
  NAND2BX1 U34 ( .AN(n144), .B(n137), .Y(n107) );
  CLKINVX1 U35 ( .A(addr[1]), .Y(n13) );
  NOR2X1 U36 ( .A(n10), .B(n3), .Y(n122) );
  NOR2X1 U37 ( .A(addr[1]), .B(n2), .Y(n132) );
  OAI22X1 U38 ( .A0(n82), .A1(n12), .B0(n5), .B1(n14), .Y(n88) );
  NAND2X1 U40 ( .A(n3), .B(n7), .Y(n123) );
  NAND4X1 U41 ( .A(n147), .B(n140), .C(n100), .D(n99), .Y(n101) );
  AOI222XL U42 ( .A0(n98), .A1(n84), .B0(n102), .B1(n130), .C0(n97), .C1(n105), 
        .Y(n99) );
  NAND3X1 U43 ( .A(n5), .B(n82), .C(n96), .Y(n100) );
  OAI221X1 U44 ( .A0(n85), .A1(n15), .B0(n82), .B1(n83), .C0(n14), .Y(n98) );
  AOI22X1 U45 ( .A0(n4), .A1(n115), .B0(addr[5]), .B1(n114), .Y(n129) );
  OAI21XL U46 ( .A0(n121), .A1(n16), .B0(n147), .Y(n115) );
  OAI21XL U48 ( .A0(n113), .A1(n84), .B0(n112), .Y(n114) );
  AOI221XL U49 ( .A0(n119), .A1(n13), .B0(n130), .B1(addr[3]), .C0(n111), .Y(
        n113) );
  OAI22XL U51 ( .A0(n12), .A1(n81), .B0(addr[3]), .B1(n10), .Y(n111) );
  OAI22XL U52 ( .A0(n85), .A1(n83), .B0(addr[1]), .B1(n82), .Y(n142) );
  AOI211X1 U53 ( .A0(n4), .A1(n135), .B0(n134), .C0(n133), .Y(n136) );
  OA21XL U54 ( .A0(n1), .A1(n3), .B0(n132), .Y(n133) );
  OAI2BB2XL U55 ( .B0(n2), .B1(n9), .A0N(n131), .A1N(n130), .Y(n134) );
  OAI22X1 U56 ( .A0(n5), .A1(n12), .B0(n84), .B1(n10), .Y(n135) );
  CLKINVX3 U57 ( .A(addr[5]), .Y(n7) );
  AOI2BB2X1 U59 ( .B0(n5), .B1(n130), .A0N(n3), .A1N(n15), .Y(n137) );
  NOR2X1 U60 ( .A(n15), .B(n2), .Y(n126) );
  AOI2BB2XL U67 ( .B0(n143), .B1(n90), .A0N(n89), .A1N(n7), .Y(n94) );
  AOI211X1 U68 ( .A0(n122), .A1(n4), .B0(n88), .C0(n87), .Y(n89) );
  OAI32X1 U69 ( .A0(n15), .A1(n85), .A2(n84), .B0(n11), .B1(n18), .Y(n87) );
  NAND3X1 U70 ( .A(n147), .B(n140), .C(n139), .Y(n141) );
  AOI32X1 U71 ( .A0(n5), .A1(n13), .A2(n4), .B0(n138), .B1(n81), .Y(n139) );
  AO22XL U72 ( .A0(n143), .A1(n2), .B0(n116), .B1(n81), .Y(n120) );
  OAI21XL U73 ( .A0(n3), .A1(n7), .B0(n123), .Y(n116) );
  CLKINVX1 U74 ( .A(n106), .Y(n8) );
  AOI32XL U75 ( .A0(n105), .A1(n81), .A2(n1), .B0(addr[1]), .B1(n125), .Y(n106) );
  OAI211X1 U76 ( .A0(n81), .A1(n140), .B0(n110), .C0(n109), .Y(dout[2]) );
  AOI222XL U77 ( .A0(n108), .A1(n7), .B0(n143), .B1(n8), .C0(n119), .C1(n107), 
        .Y(n109) );
  AOI2BB2XL U78 ( .B0(addr[5]), .B1(n101), .A0N(n84), .A1N(n112), .Y(n110) );
  OAI211X1 U79 ( .A0(n2), .A1(n147), .B0(n146), .C0(n145), .Y(dout[4]) );
  AOI222XL U80 ( .A0(n144), .A1(n85), .B0(n143), .B1(n142), .C0(n141), .C1(n7), 
        .Y(n145) );
  OA22X1 U81 ( .A0(n17), .A1(n137), .B0(n136), .B1(n7), .Y(n146) );
  NAND3X1 U82 ( .A(n129), .B(n128), .C(n127), .Y(dout[3]) );
  AOI32XL U83 ( .A0(n120), .A1(n85), .A2(addr[1]), .B0(n119), .B1(n118), .Y(
        n128) );
  AOI222XL U84 ( .A0(n144), .A1(n81), .B0(n126), .B1(n6), .C0(n125), .C1(n124), 
        .Y(n127) );
  NAND3BX1 U85 ( .AN(n95), .B(n94), .C(n93), .Y(dout[1]) );
  OAI222X1 U86 ( .A0(n140), .A1(n4), .B0(n112), .B1(n84), .C0(n10), .C1(n91), 
        .Y(n95) );
  AOI32XL U87 ( .A0(addr[1]), .A1(n7), .A2(n125), .B0(n130), .B1(n92), .Y(n93)
         );
  CLKINVX3 U88 ( .A(addr[6]), .Y(n83) );
  CLKINVX3 U89 ( .A(n5), .Y(n84) );
endmodule


module sbox7_4 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148;

  OAI222X4 U19 ( .A0(n20), .A1(n129), .B0(n4), .B1(n16), .C0(addr[1]), .C1(n8), 
        .Y(n122) );
  OAI33X4 U33 ( .A0(addr[1]), .A1(n4), .A2(n5), .B0(n17), .B1(n6), .B2(n14), 
        .Y(n97) );
  NOR2X2 U44 ( .A(n84), .B(n4), .Y(n116) );
  NOR2X2 U48 ( .A(addr[1]), .B(addr[6]), .Y(n136) );
  NOR2X2 U51 ( .A(n87), .B(n84), .Y(n125) );
  NOR2X2 U52 ( .A(n17), .B(addr[3]), .Y(n131) );
  NOR2X2 U58 ( .A(n93), .B(n124), .Y(n142) );
  NOR2X2 U60 ( .A(n86), .B(addr[1]), .Y(n93) );
  NOR2X2 U62 ( .A(n12), .B(n3), .Y(n137) );
  NOR2X2 U65 ( .A(n86), .B(n18), .Y(n140) );
  NAND2X1 U1 ( .A(n3), .B(n4), .Y(n119) );
  CLKBUFX3 U2 ( .A(addr[4]), .Y(n4) );
  CLKINVX1 U3 ( .A(n12), .Y(n1) );
  CLKINVX1 U4 ( .A(n6), .Y(n2) );
  CLKBUFX3 U5 ( .A(addr[2]), .Y(n5) );
  OAI31X1 U6 ( .A0(n84), .A1(n12), .A2(n18), .B0(n117), .Y(n121) );
  NOR2X4 U7 ( .A(n18), .B(addr[6]), .Y(n124) );
  OAI22X1 U8 ( .A0(addr[1]), .A1(n8), .B0(n5), .B1(n113), .Y(n100) );
  OAI22X1 U9 ( .A0(n4), .A1(n87), .B0(addr[3]), .B1(n11), .Y(n103) );
  AOI211XL U10 ( .A0(n5), .A1(n15), .B0(n131), .C0(n130), .Y(n132) );
  NOR3XL U11 ( .A(n20), .B(addr[3]), .C(n2), .Y(n130) );
  OAI21XL U12 ( .A0(n3), .A1(n1), .B0(n119), .Y(n89) );
  BUFX4 U13 ( .A(addr[5]), .Y(n3) );
  AOI221XL U14 ( .A0(n140), .A1(n89), .B0(n109), .B1(n15), .C0(n88), .Y(n96)
         );
  CLKINVX1 U15 ( .A(n140), .Y(n17) );
  OAI2BB2XL U16 ( .B0(n142), .B1(n11), .A0N(n141), .A1N(n140), .Y(n143) );
  CLKINVX1 U17 ( .A(n125), .Y(n83) );
  CLKINVX1 U18 ( .A(n142), .Y(n15) );
  NAND2X1 U20 ( .A(n83), .B(n85), .Y(n105) );
  CLKINVX1 U21 ( .A(n123), .Y(n7) );
  CLKINVX1 U22 ( .A(n109), .Y(n10) );
  NAND2X1 U23 ( .A(n124), .B(n84), .Y(n113) );
  CLKINVX1 U24 ( .A(n137), .Y(n11) );
  NOR2X1 U25 ( .A(n11), .B(n84), .Y(n109) );
  CLKINVX1 U26 ( .A(n136), .Y(n20) );
  OAI22XL U27 ( .A0(n137), .A1(n16), .B0(n18), .B1(n10), .Y(n146) );
  OAI21X1 U28 ( .A0(n12), .A1(n83), .B0(n129), .Y(n141) );
  NAND2X1 U29 ( .A(n116), .B(n87), .Y(n129) );
  CLKINVX1 U30 ( .A(n93), .Y(n19) );
  OAI21XL U31 ( .A0(n119), .A1(n19), .B0(n118), .Y(n120) );
  OAI21XL U32 ( .A0(n125), .A1(n137), .B0(n124), .Y(n118) );
  NOR2X1 U34 ( .A(n87), .B(n8), .Y(n123) );
  CLKINVX1 U35 ( .A(n145), .Y(n8) );
  OAI22XL U36 ( .A0(n137), .A1(n113), .B0(n86), .B1(n7), .Y(n88) );
  CLKINVX1 U37 ( .A(n116), .Y(n14) );
  CLKINVX1 U38 ( .A(n131), .Y(n16) );
  CLKINVX1 U39 ( .A(n134), .Y(n85) );
  NOR2XL U40 ( .A(n125), .B(n12), .Y(n110) );
  CLKINVX1 U41 ( .A(n119), .Y(n13) );
  CLKINVX1 U42 ( .A(n103), .Y(n9) );
  OA21XL U43 ( .A0(n21), .A1(n19), .B0(n117), .Y(n102) );
  CLKINVX1 U45 ( .A(n105), .Y(n21) );
  OAI2BB1XL U46 ( .A0N(n103), .A1N(n124), .B0(n102), .Y(n104) );
  OAI22X1 U47 ( .A0(n87), .A1(n14), .B0(n4), .B1(n85), .Y(n112) );
  NOR4X1 U49 ( .A(n4), .B(addr[3]), .C(n18), .D(n6), .Y(n99) );
  XNOR2X1 U50 ( .A(addr[6]), .B(n5), .Y(n101) );
  AOI211X1 U53 ( .A0(n116), .A1(addr[6]), .B0(n115), .C0(n114), .Y(n128) );
  OAI222X1 U54 ( .A0(n111), .A1(n17), .B0(n110), .B1(n19), .C0(n20), .C1(n10), 
        .Y(n115) );
  OAI2BB2XL U55 ( .B0(n13), .B1(n113), .A0N(n18), .A1N(n112), .Y(n114) );
  OA21XL U56 ( .A0(n84), .A1(n3), .B0(n7), .Y(n111) );
  NAND2X1 U57 ( .A(n5), .B(n136), .Y(n133) );
  CLKINVX1 U59 ( .A(addr[6]), .Y(n86) );
  AOI211X1 U61 ( .A0(n131), .A1(n3), .B0(n92), .C0(n91), .Y(n95) );
  OAI221X1 U63 ( .A0(n18), .A1(n8), .B0(n17), .B1(n11), .C0(n102), .Y(n92) );
  OAI31X1 U64 ( .A0(n84), .A1(n12), .A2(n20), .B0(n90), .Y(n91) );
  AO21XL U66 ( .A0(n119), .A1(n129), .B0(addr[6]), .Y(n90) );
  NOR2X1 U67 ( .A(n12), .B(addr[3]), .Y(n145) );
  AOI21XL U68 ( .A0(addr[3]), .A1(n98), .B0(n97), .Y(n108) );
  OAI2BB1XL U69 ( .A0N(n6), .A1N(n124), .B0(n133), .Y(n98) );
  NAND3X1 U70 ( .A(n136), .B(n84), .C(n3), .Y(n117) );
  NOR2X1 U71 ( .A(addr[3]), .B(n3), .Y(n134) );
  OAI21X1 U72 ( .A0(n5), .A1(n142), .B0(n133), .Y(n138) );
  OAI22XL U73 ( .A0(n142), .A1(n14), .B0(n1), .B1(n132), .Y(n135) );
  AO21X1 U74 ( .A0(n139), .A1(n87), .B0(n138), .Y(n144) );
  OAI21XL U75 ( .A0(n2), .A1(n18), .B0(n19), .Y(n139) );
  OAI221X1 U76 ( .A0(n96), .A1(n6), .B0(n5), .B1(n95), .C0(n94), .Y(dout[1])
         );
  AOI2BB2X1 U77 ( .B0(n93), .B1(n112), .A0N(n133), .A1N(n9), .Y(n94) );
  OAI211X1 U78 ( .A0(n128), .A1(n6), .B0(n127), .C0(n126), .Y(dout[3]) );
  AOI32XL U79 ( .A0(n125), .A1(n1), .A2(n124), .B0(n123), .B1(n136), .Y(n126)
         );
  OAI31X1 U80 ( .A0(n122), .A1(n121), .A2(n120), .B0(n6), .Y(n127) );
  OAI221X1 U81 ( .A0(n3), .A1(n108), .B0(n107), .B1(n87), .C0(n106), .Y(
        dout[2]) );
  AOI32XL U82 ( .A0(n105), .A1(n6), .A2(n140), .B0(n2), .B1(n104), .Y(n106) );
  AOI211X1 U83 ( .A0(n101), .A1(n4), .B0(n100), .C0(n99), .Y(n107) );
  NAND2X1 U84 ( .A(n148), .B(n147), .Y(dout[4]) );
  AOI222XL U85 ( .A0(n136), .A1(n141), .B0(n3), .B1(n135), .C0(n134), .C1(n138), .Y(n148) );
  AOI222XL U86 ( .A0(n5), .A1(n146), .B0(n145), .B1(n144), .C0(n143), .C1(n6), 
        .Y(n147) );
  CLKINVX3 U87 ( .A(n5), .Y(n6) );
  CLKINVX3 U88 ( .A(n4), .Y(n12) );
  CLKINVX3 U89 ( .A(addr[1]), .Y(n18) );
  CLKINVX3 U90 ( .A(addr[3]), .Y(n84) );
  CLKINVX3 U91 ( .A(n3), .Y(n87) );
endmodule


module sbox8_4 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132;

  NAND2X2 U41 ( .A(addr[6]), .B(n9), .Y(n131) );
  NAND2X2 U48 ( .A(addr[4]), .B(n6), .Y(n123) );
  NAND2X2 U49 ( .A(n2), .B(n74), .Y(n87) );
  NAND2X2 U50 ( .A(addr[1]), .B(n16), .Y(n124) );
  NAND2X2 U54 ( .A(addr[2]), .B(n14), .Y(n116) );
  NAND2X2 U60 ( .A(addr[6]), .B(addr[1]), .Y(n105) );
  NAND2X2 U61 ( .A(n9), .B(n16), .Y(n108) );
  OAI32X1 U1 ( .A0(n16), .A1(addr[4]), .A2(n92), .B0(n115), .B1(n108), .Y(n96)
         );
  OAI31X1 U2 ( .A0(n123), .A1(addr[6]), .A2(n116), .B0(n109), .Y(n110) );
  OAI221X1 U3 ( .A0(n105), .A1(n87), .B0(addr[4]), .B1(n108), .C0(n86), .Y(n90) );
  NAND2X4 U4 ( .A(addr[4]), .B(n2), .Y(n115) );
  AOI222X1 U5 ( .A0(n88), .A1(addr[2]), .B0(n74), .B1(n15), .C0(n75), .C1(n92), 
        .Y(n114) );
  OAI222X1 U6 ( .A0(addr[2]), .A1(n126), .B0(n6), .B1(n125), .C0(n124), .C1(
        n123), .Y(n127) );
  AOI32XL U7 ( .A0(n12), .A1(n13), .A2(n2), .B0(n8), .B1(n117), .Y(n130) );
  OA21XL U8 ( .A0(n75), .A1(n14), .B0(n121), .Y(n78) );
  INVXL U9 ( .A(n119), .Y(n3) );
  INVX3 U10 ( .A(n2), .Y(n6) );
  BUFX4 U11 ( .A(addr[3]), .Y(n2) );
  CLKBUFX3 U12 ( .A(addr[5]), .Y(n1) );
  CLKINVX1 U13 ( .A(n108), .Y(n8) );
  CLKINVX1 U14 ( .A(n107), .Y(n4) );
  CLKINVX1 U15 ( .A(n93), .Y(n5) );
  NAND2X1 U16 ( .A(n6), .B(n74), .Y(n93) );
  NAND2X1 U17 ( .A(n75), .B(n14), .Y(n121) );
  OAI21XL U18 ( .A0(n115), .A1(n14), .B0(n107), .Y(n77) );
  OAI21X1 U19 ( .A0(n74), .A1(n14), .B0(n123), .Y(n88) );
  OAI31XL U20 ( .A0(n115), .A1(n9), .A2(n116), .B0(n118), .Y(n94) );
  CLKINVX1 U21 ( .A(n131), .Y(n7) );
  NAND2X1 U22 ( .A(n13), .B(n6), .Y(n107) );
  OAI22XL U23 ( .A0(n116), .A1(n123), .B0(n13), .B1(n115), .Y(n117) );
  OAI22XL U24 ( .A0(n123), .A1(n108), .B0(n131), .B1(n93), .Y(n95) );
  OAI2BB2XL U25 ( .B0(n115), .B1(n131), .A0N(n88), .A1N(n11), .Y(n89) );
  AOI211XL U26 ( .A0(n108), .A1(n105), .B0(n74), .C0(n121), .Y(n85) );
  CLKINVX1 U27 ( .A(n124), .Y(n12) );
  OAI22XL U28 ( .A0(n13), .A1(n123), .B0(n78), .B1(n87), .Y(n81) );
  NAND2BX2 U29 ( .AN(n78), .B(n6), .Y(n120) );
  NAND2XL U30 ( .A(n115), .B(n93), .Y(n104) );
  OAI2BB2XL U31 ( .B0(n106), .B1(n105), .A0N(n104), .A1N(n12), .Y(n111) );
  NOR2BXL U32 ( .AN(n123), .B(n103), .Y(n106) );
  NAND3X1 U33 ( .A(n104), .B(n9), .C(n13), .Y(n84) );
  AO21X1 U34 ( .A0(n13), .A1(n11), .B0(n101), .Y(n102) );
  OAI33X1 U35 ( .A0(n16), .A1(n6), .A2(n100), .B0(n75), .B1(n103), .B2(n124), 
        .Y(n101) );
  OA22XL U36 ( .A0(n107), .A1(n131), .B0(n120), .B1(n124), .Y(n98) );
  CLKINVX1 U37 ( .A(n125), .Y(n10) );
  OAI21XL U38 ( .A0(n12), .A1(n7), .B0(addr[4]), .Y(n86) );
  NAND2X1 U39 ( .A(n1), .B(n75), .Y(n100) );
  OAI221X1 U40 ( .A0(n124), .A1(n121), .B0(addr[1]), .B1(n120), .C0(n3), .Y(
        n128) );
  OAI31XL U42 ( .A0(n75), .A1(n9), .A2(n6), .B0(n118), .Y(n119) );
  NAND2X1 U43 ( .A(n11), .B(addr[2]), .Y(n125) );
  NAND4XL U44 ( .A(n7), .B(n1), .C(n2), .D(addr[2]), .Y(n109) );
  NAND3X1 U45 ( .A(n13), .B(n16), .C(n2), .Y(n118) );
  OAI21XL U46 ( .A0(n1), .A1(n87), .B0(n114), .Y(n76) );
  OAI22XL U47 ( .A0(n108), .A1(n120), .B0(n79), .B1(n100), .Y(n80) );
  AOI221XL U51 ( .A0(n7), .A1(n6), .B0(n11), .B1(n2), .C0(n91), .Y(n79) );
  NOR2X1 U52 ( .A(n1), .B(n2), .Y(n103) );
  NOR2X1 U53 ( .A(n87), .B(addr[6]), .Y(n91) );
  NOR2X1 U55 ( .A(n6), .B(n1), .Y(n92) );
  CLKINVX1 U56 ( .A(n100), .Y(n15) );
  OA21XL U57 ( .A0(n1), .A1(n115), .B0(n120), .Y(n132) );
  AOI221XL U58 ( .A0(n8), .A1(n2), .B0(n11), .B1(addr[4]), .C0(n122), .Y(n126)
         );
  OAI22XL U59 ( .A0(n2), .A1(n9), .B0(addr[4]), .B1(n131), .Y(n122) );
  OAI211X1 U62 ( .A0(addr[2]), .A1(n99), .B0(n98), .C0(n97), .Y(dout[2]) );
  AOI221XL U63 ( .A0(addr[2]), .A1(n96), .B0(n1), .B1(n95), .C0(n94), .Y(n97)
         );
  AOI221XL U64 ( .A0(n91), .A1(n1), .B0(n90), .B1(n14), .C0(n89), .Y(n99) );
  OAI211X1 U65 ( .A0(n132), .A1(n131), .B0(n130), .C0(n129), .Y(dout[4]) );
  AOI222XL U66 ( .A0(n128), .A1(n74), .B0(n1), .B1(n127), .C0(n4), .C1(n11), 
        .Y(n129) );
  OAI211X1 U67 ( .A0(addr[1]), .A1(n114), .B0(n113), .C0(n112), .Y(dout[3]) );
  AOI221XL U68 ( .A0(n111), .A1(n75), .B0(n4), .B1(n8), .C0(n110), .Y(n112) );
  AOI2BB2XL U69 ( .B0(n102), .B1(n74), .A0N(n115), .A1N(n125), .Y(n113) );
  NAND4BX1 U70 ( .AN(n85), .B(n84), .C(n83), .D(n82), .Y(dout[1]) );
  AOI221XL U71 ( .A0(n7), .A1(n81), .B0(n5), .B1(n10), .C0(n80), .Y(n82) );
  AOI22X1 U72 ( .A0(n11), .A1(n77), .B0(n12), .B1(n76), .Y(n83) );
  CLKINVX3 U73 ( .A(addr[1]), .Y(n9) );
  CLKINVX3 U74 ( .A(n105), .Y(n11) );
  CLKINVX3 U75 ( .A(n116), .Y(n13) );
  CLKINVX3 U76 ( .A(n1), .Y(n14) );
  CLKINVX3 U77 ( .A(addr[6]), .Y(n16) );
  CLKINVX3 U78 ( .A(addr[4]), .Y(n74) );
  CLKINVX3 U79 ( .A(addr[2]), .Y(n75) );
endmodule


module crp_4 ( P, R, K_sub );
  output [1:32] P;
  input [1:32] R;
  input [1:48] K_sub;
  wire   n1;
  wire   [1:48] X;

  sbox1_4 u0 ( .addr(X[1:6]), .dout({P[9], P[17], P[23], P[31]}) );
  sbox2_4 u1 ( .addr({X[7], n1, X[9:12]}), .dout({P[13], P[28], P[2], P[18]})
         );
  sbox3_4 u2 ( .addr(X[13:18]), .dout({P[24], P[16], P[30], P[6]}) );
  sbox4_4 u3 ( .addr(X[19:24]), .dout({P[26], P[20], P[10], P[1]}) );
  sbox5_4 u4 ( .addr(X[25:30]), .dout({P[8], P[14], P[25], P[3]}) );
  sbox6_4 u5 ( .addr(X[31:36]), .dout({P[4], P[29], P[11], P[19]}) );
  sbox7_4 u6 ( .addr(X[37:42]), .dout({P[32], P[12], P[22], P[7]}) );
  sbox8_4 u7 ( .addr(X[43:48]), .dout({P[5], P[27], P[15], P[21]}) );
  XOR2X1 U1 ( .A(R[1]), .B(K_sub[2]), .Y(X[2]) );
  CLKXOR2X4 U2 ( .A(R[10]), .B(K_sub[15]), .Y(X[15]) );
  CLKXOR2X4 U3 ( .A(R[29]), .B(K_sub[42]), .Y(X[42]) );
  CLKXOR2X4 U4 ( .A(R[5]), .B(K_sub[6]), .Y(X[6]) );
  CLKXOR2X4 U5 ( .A(R[8]), .B(K_sub[11]), .Y(X[11]) );
  CLKXOR2X4 U6 ( .A(R[16]), .B(K_sub[25]), .Y(X[25]) );
  CLKXOR2X4 U7 ( .A(R[20]), .B(K_sub[31]), .Y(X[31]) );
  CLKXOR2X4 U8 ( .A(R[16]), .B(K_sub[23]), .Y(X[23]) );
  XNOR2X1 U9 ( .A(R[5]), .B(K_sub[8]), .Y(X[8]) );
  INVX3 U10 ( .A(X[8]), .Y(n1) );
  CLKXOR2X4 U11 ( .A(R[31]), .B(K_sub[46]), .Y(X[46]) );
  CLKXOR2X4 U12 ( .A(R[22]), .B(K_sub[33]), .Y(X[33]) );
  CLKXOR2X4 U13 ( .A(R[29]), .B(K_sub[44]), .Y(X[44]) );
  CLKXOR2X4 U14 ( .A(R[12]), .B(K_sub[19]), .Y(X[19]) );
  CLKXOR2X4 U15 ( .A(R[26]), .B(K_sub[39]), .Y(X[39]) );
  CLKXOR2X4 U16 ( .A(R[20]), .B(K_sub[29]), .Y(X[29]) );
  CLKXOR2X2 U17 ( .A(R[4]), .B(K_sub[5]), .Y(X[5]) );
  CLKXOR2X2 U18 ( .A(R[15]), .B(K_sub[22]), .Y(X[22]) );
  CLKXOR2X2 U19 ( .A(R[24]), .B(K_sub[35]), .Y(X[35]) );
  CLKXOR2X2 U20 ( .A(R[21]), .B(K_sub[30]), .Y(X[30]) );
  CLKXOR2X2 U21 ( .A(R[12]), .B(K_sub[17]), .Y(X[17]) );
  CLKXOR2X2 U22 ( .A(R[32]), .B(K_sub[1]), .Y(X[1]) );
  CLKXOR2X2 U23 ( .A(R[13]), .B(K_sub[20]), .Y(X[20]) );
  CLKXOR2X2 U24 ( .A(R[18]), .B(K_sub[27]), .Y(X[27]) );
  CLKXOR2X2 U25 ( .A(R[8]), .B(K_sub[13]), .Y(X[13]) );
  CLKXOR2X2 U26 ( .A(R[4]), .B(K_sub[7]), .Y(X[7]) );
  CLKXOR2X2 U27 ( .A(R[24]), .B(K_sub[37]), .Y(X[37]) );
  CLKXOR2X2 U28 ( .A(R[28]), .B(K_sub[43]), .Y(X[43]) );
  CLKXOR2X2 U29 ( .A(R[1]), .B(K_sub[48]), .Y(X[48]) );
  CLKXOR2X2 U30 ( .A(R[17]), .B(K_sub[24]), .Y(X[24]) );
  CLKXOR2X2 U31 ( .A(R[9]), .B(K_sub[12]), .Y(X[12]) );
  CLKXOR2X2 U32 ( .A(R[13]), .B(K_sub[18]), .Y(X[18]) );
  CLKXOR2X2 U33 ( .A(R[25]), .B(K_sub[36]), .Y(X[36]) );
  XOR2X1 U34 ( .A(R[23]), .B(K_sub[34]), .Y(X[34]) );
  XOR2X1 U35 ( .A(R[9]), .B(K_sub[14]), .Y(X[14]) );
  XOR2X1 U36 ( .A(R[30]), .B(K_sub[45]), .Y(X[45]) );
  XOR2X1 U37 ( .A(R[21]), .B(K_sub[32]), .Y(X[32]) );
  XOR2X1 U38 ( .A(R[25]), .B(K_sub[38]), .Y(X[38]) );
  XOR2X1 U39 ( .A(R[27]), .B(K_sub[40]), .Y(X[40]) );
  XOR2X1 U40 ( .A(R[3]), .B(K_sub[4]), .Y(X[4]) );
  XOR2X1 U41 ( .A(R[11]), .B(K_sub[16]), .Y(X[16]) );
  XOR2X1 U42 ( .A(R[7]), .B(K_sub[10]), .Y(X[10]) );
  XOR2X1 U43 ( .A(R[14]), .B(K_sub[21]), .Y(X[21]) );
  XOR2X1 U44 ( .A(R[6]), .B(K_sub[9]), .Y(X[9]) );
  XOR2X1 U45 ( .A(R[2]), .B(K_sub[3]), .Y(X[3]) );
  XOR2X1 U46 ( .A(R[28]), .B(K_sub[41]), .Y(X[41]) );
  XOR2X1 U47 ( .A(R[17]), .B(K_sub[26]), .Y(X[26]) );
  XOR2X1 U48 ( .A(R[32]), .B(K_sub[47]), .Y(X[47]) );
  XOR2X1 U49 ( .A(R[19]), .B(K_sub[28]), .Y(X[28]) );
endmodule


module sbox1_3 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127;

  OAI222X4 U13 ( .A0(addr[5]), .A1(n101), .B0(n1), .B1(n100), .C0(n99), .C1(n9), .Y(dout[3]) );
  OAI21X2 U42 ( .A0(n4), .A1(n112), .B0(n106), .Y(n123) );
  NAND2X2 U44 ( .A(addr[6]), .B(n69), .Y(n115) );
  NAND2X2 U48 ( .A(addr[1]), .B(n72), .Y(n114) );
  OAI22X2 U49 ( .A0(n11), .A1(n10), .B0(addr[5]), .B1(n120), .Y(n85) );
  NAND2X2 U50 ( .A(n3), .B(n11), .Y(n120) );
  NOR2X2 U51 ( .A(n11), .B(n3), .Y(n124) );
  NOR2X2 U56 ( .A(n109), .B(n3), .Y(n93) );
  NAND2X2 U57 ( .A(addr[1]), .B(addr[6]), .Y(n109) );
  NAND2X2 U59 ( .A(n69), .B(n72), .Y(n112) );
  NOR2X1 U1 ( .A(n114), .B(n120), .Y(n104) );
  AOI221X4 U2 ( .A0(n13), .A1(n90), .B0(n4), .B1(n93), .C0(n102), .Y(n79) );
  NOR3X1 U3 ( .A(n2), .B(addr[6]), .C(n9), .Y(n102) );
  BUFX4 U4 ( .A(addr[4]), .Y(n2) );
  CLKBUFX3 U5 ( .A(addr[2]), .Y(n1) );
  OAI32X1 U6 ( .A0(n112), .A1(n2), .A2(n4), .B0(n115), .B1(n113), .Y(n80) );
  NOR2BXL U7 ( .AN(n118), .B(n1), .Y(n122) );
  CLKBUFX3 U8 ( .A(addr[2]), .Y(n4) );
  OAI221X4 U9 ( .A0(n88), .A1(n10), .B0(addr[5]), .B1(n87), .C0(n86), .Y(
        dout[2]) );
  OAI221X4 U10 ( .A0(addr[5]), .A1(n127), .B0(n126), .B1(n10), .C0(n125), .Y(
        dout[4]) );
  OA21XL U11 ( .A0(n95), .A1(n115), .B0(n107), .Y(n119) );
  AOI222XL U12 ( .A0(n13), .A1(n1), .B0(n2), .B1(n110), .C0(n70), .C1(n9), .Y(
        n111) );
  AOI2BB2X1 U14 ( .B0(n2), .B1(n70), .A0N(addr[4]), .A1N(n115), .Y(n91) );
  BUFX4 U15 ( .A(addr[3]), .Y(n3) );
  CLKINVX1 U16 ( .A(n112), .Y(n13) );
  CLKINVX1 U17 ( .A(n113), .Y(n5) );
  NAND2BX1 U18 ( .AN(n104), .B(n119), .Y(n84) );
  CLKXOR2X2 U19 ( .A(n6), .B(n9), .Y(n90) );
  NOR2X1 U20 ( .A(n11), .B(n6), .Y(n118) );
  OAI21XL U21 ( .A0(n6), .A1(n114), .B0(n91), .Y(n92) );
  NAND2X1 U22 ( .A(n93), .B(n11), .Y(n107) );
  NAND2X1 U23 ( .A(n9), .B(n6), .Y(n113) );
  OAI211X1 U24 ( .A0(n11), .A1(n114), .B0(n108), .C0(n107), .Y(n89) );
  CLKINVX1 U25 ( .A(n109), .Y(n70) );
  NAND2X1 U26 ( .A(n124), .B(n12), .Y(n108) );
  CLKINVX1 U27 ( .A(n114), .Y(n71) );
  CLKINVX1 U28 ( .A(n115), .Y(n12) );
  CLKINVX1 U29 ( .A(n95), .Y(n8) );
  AO22X1 U30 ( .A0(n90), .A1(n12), .B0(n6), .B1(n123), .Y(n76) );
  OAI31X1 U31 ( .A0(n9), .A1(n3), .A2(n69), .B0(n103), .Y(n105) );
  AOI31XL U32 ( .A0(n69), .A1(n9), .A2(n2), .B0(n102), .Y(n103) );
  CLKINVX1 U33 ( .A(addr[6]), .Y(n72) );
  AOI211X1 U34 ( .A0(n7), .A1(n4), .B0(n117), .C0(n116), .Y(n126) );
  CLKINVX1 U35 ( .A(n108), .Y(n7) );
  AOI211X1 U36 ( .A0(n115), .A1(n114), .B0(n113), .C0(n2), .Y(n116) );
  OAI22X1 U37 ( .A0(n120), .A1(n112), .B0(n111), .B1(n6), .Y(n117) );
  AOI211X1 U38 ( .A0(n70), .A1(n118), .B0(n81), .C0(n80), .Y(n88) );
  OAI22X1 U39 ( .A0(n91), .A1(n9), .B0(n3), .B1(n106), .Y(n81) );
  CLKINVX3 U40 ( .A(addr[5]), .Y(n10) );
  NAND2X1 U41 ( .A(n3), .B(n10), .Y(n95) );
  NAND2X1 U43 ( .A(n71), .B(n1), .Y(n106) );
  XOR2X1 U45 ( .A(n82), .B(n2), .Y(n83) );
  NAND2X1 U46 ( .A(n1), .B(n3), .Y(n82) );
  OAI22XL U47 ( .A0(n3), .A1(n69), .B0(n6), .B1(n112), .Y(n94) );
  AOI211XL U52 ( .A0(n98), .A1(n6), .B0(n97), .C0(n104), .Y(n99) );
  OAI22XL U53 ( .A0(n96), .A1(n11), .B0(n95), .B1(n109), .Y(n97) );
  OAI22XL U54 ( .A0(n72), .A1(n10), .B0(n2), .B1(addr[1]), .Y(n98) );
  AOI221XL U55 ( .A0(n8), .A1(addr[6]), .B0(addr[5]), .B1(n94), .C0(n93), .Y(
        n96) );
  OAI21XL U58 ( .A0(addr[1]), .A1(n120), .B0(n119), .Y(n121) );
  AOI221XL U60 ( .A0(n13), .A1(n118), .B0(n93), .B1(n10), .C0(n75), .Y(n78) );
  OAI31X1 U61 ( .A0(n10), .A1(n2), .A2(n74), .B0(n73), .Y(n75) );
  OA21XL U62 ( .A0(n3), .A1(n72), .B0(n109), .Y(n74) );
  OAI21XL U63 ( .A0(n124), .A1(n85), .B0(n71), .Y(n73) );
  OAI21XL U64 ( .A0(n1), .A1(n69), .B0(n109), .Y(n110) );
  INVX4 U65 ( .A(n4), .Y(n9) );
  AOI222XL U66 ( .A0(n124), .A1(n123), .B0(n122), .B1(addr[6]), .C0(n1), .C1(
        n121), .Y(n125) );
  NOR4BBX1 U67 ( .AN(n107), .BN(n106), .C(n105), .D(n104), .Y(n127) );
  AOI222XL U68 ( .A0(n13), .A1(n90), .B0(n89), .B1(n9), .C0(n123), .C1(n11), 
        .Y(n101) );
  AOI2BB2XL U69 ( .B0(addr[5]), .B1(n92), .A0N(n120), .A1N(addr[1]), .Y(n100)
         );
  AOI32X1 U70 ( .A0(n4), .A1(n85), .A2(n13), .B0(n84), .B1(n9), .Y(n86) );
  AOI222XL U71 ( .A0(n124), .A1(n69), .B0(n83), .B1(addr[1]), .C0(n5), .C1(n72), .Y(n87) );
  OAI221X1 U72 ( .A0(n79), .A1(n10), .B0(n4), .B1(n78), .C0(n77), .Y(dout[1])
         );
  AOI32XL U73 ( .A0(addr[6]), .A1(n85), .A2(n1), .B0(n76), .B1(n10), .Y(n77)
         );
  CLKINVX3 U74 ( .A(n3), .Y(n6) );
  CLKINVX3 U75 ( .A(n2), .Y(n11) );
  CLKINVX3 U76 ( .A(addr[1]), .Y(n69) );
endmodule


module sbox2_3 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147;

  NAND2X2 U55 ( .A(n2), .B(n16), .Y(n136) );
  NAND2X2 U57 ( .A(addr[2]), .B(n83), .Y(n104) );
  NAND2X2 U60 ( .A(addr[5]), .B(addr[2]), .Y(n132) );
  NOR2X2 U61 ( .A(n7), .B(n4), .Y(n101) );
  NAND2X2 U62 ( .A(n6), .B(n9), .Y(n146) );
  NAND2X2 U63 ( .A(n3), .B(n11), .Y(n124) );
  NAND2X2 U64 ( .A(addr[6]), .B(n6), .Y(n122) );
  NAND2X2 U67 ( .A(n3), .B(n2), .Y(n133) );
  AOI222XL U1 ( .A0(n15), .A1(n8), .B0(n88), .B1(n11), .C0(n140), .C1(n4), .Y(
        n89) );
  CLKINVX1 U2 ( .A(n121), .Y(n7) );
  OAI211X4 U3 ( .A0(n147), .A1(n146), .B0(n145), .C0(n144), .Y(dout[4]) );
  NOR2X1 U4 ( .A(n104), .B(n2), .Y(n141) );
  NOR2X1 U5 ( .A(n124), .B(n2), .Y(n140) );
  CLKBUFX4 U6 ( .A(addr[4]), .Y(n2) );
  CLKINVX1 U7 ( .A(addr[5]), .Y(n1) );
  INVX3 U8 ( .A(addr[5]), .Y(n83) );
  NAND3XL U9 ( .A(n98), .B(n97), .C(n96), .Y(dout[1]) );
  NAND2X1 U10 ( .A(addr[1]), .B(addr[6]), .Y(n121) );
  CLKINVX2 U11 ( .A(addr[1]), .Y(n6) );
  OAI221X1 U12 ( .A0(addr[1]), .A1(n136), .B0(n133), .B1(n6), .C0(n87), .Y(n95) );
  NAND2X4 U13 ( .A(addr[1]), .B(n9), .Y(n114) );
  INVX3 U14 ( .A(addr[6]), .Y(n9) );
  NAND2XL U15 ( .A(n102), .B(n16), .Y(n109) );
  AOI211XL U16 ( .A0(n12), .A1(n95), .B0(n94), .C0(n93), .Y(n96) );
  AOI2BB2X1 U17 ( .B0(n83), .B1(n10), .A0N(n104), .A1N(n136), .Y(n117) );
  NOR3BXL U18 ( .AN(n135), .B(n134), .C(n15), .Y(n147) );
  BUFX4 U19 ( .A(addr[3]), .Y(n3) );
  NAND2X1 U20 ( .A(n15), .B(n7), .Y(n113) );
  CLKINVX1 U21 ( .A(n146), .Y(n4) );
  CLKINVX1 U22 ( .A(n115), .Y(n15) );
  CLKINVX1 U23 ( .A(n122), .Y(n5) );
  OAI31X1 U24 ( .A0(n124), .A1(n9), .A2(n83), .B0(n123), .Y(n128) );
  OAI21XL U25 ( .A0(n83), .A1(n6), .B0(n140), .Y(n123) );
  OAI22X1 U26 ( .A0(n122), .A1(n124), .B0(n101), .B1(n132), .Y(n84) );
  INVX1 U27 ( .A(n114), .Y(n8) );
  OAI22X1 U28 ( .A0(n122), .A1(n16), .B0(n82), .B1(n121), .Y(n129) );
  NAND3X1 U29 ( .A(n82), .B(n83), .C(n6), .Y(n111) );
  NAND2X1 U30 ( .A(n16), .B(n82), .Y(n115) );
  OAI21XL U31 ( .A0(n11), .A1(n133), .B0(n135), .Y(n85) );
  OAI22XL U32 ( .A0(n117), .A1(n146), .B0(n116), .B1(n132), .Y(n118) );
  AOI222XL U33 ( .A0(n8), .A1(n115), .B0(n81), .B1(n9), .C0(n15), .C1(n4), .Y(
        n116) );
  CLKINVX1 U34 ( .A(n104), .Y(n13) );
  OAI2BB2XL U35 ( .B0(n114), .B1(n135), .A0N(n126), .A1N(n81), .Y(n106) );
  OAI21XL U36 ( .A0(n112), .A1(n114), .B0(n111), .Y(n120) );
  OAI21XL U37 ( .A0(n133), .A1(n114), .B0(n113), .Y(n119) );
  CLKINVX1 U38 ( .A(n124), .Y(n10) );
  CLKINVX1 U39 ( .A(n136), .Y(n14) );
  CLKINVX1 U40 ( .A(n133), .Y(n81) );
  CLKINVX1 U41 ( .A(n132), .Y(n12) );
  AOI2BB1X1 U42 ( .A0N(n126), .A1N(n125), .B0(n136), .Y(n127) );
  OAI22XL U43 ( .A0(n104), .A1(n114), .B0(n101), .B1(n132), .Y(n102) );
  AO21XL U44 ( .A0(n11), .A1(n14), .B0(n141), .Y(n86) );
  AO21X1 U45 ( .A0(n16), .A1(n13), .B0(n140), .Y(n142) );
  NAND3X1 U46 ( .A(n11), .B(n82), .C(addr[5]), .Y(n135) );
  OAI22X1 U47 ( .A0(addr[5]), .A1(n121), .B0(n122), .B1(n83), .Y(n126) );
  AOI2BB1X1 U48 ( .A0N(n3), .A1N(n1), .B0(n14), .Y(n112) );
  NOR3X1 U49 ( .A(addr[1]), .B(addr[2]), .C(n83), .Y(n125) );
  AOI2BB1XL U50 ( .A0N(n92), .A1N(n91), .B0(addr[5]), .Y(n93) );
  OAI22XL U51 ( .A0(n117), .A1(n114), .B0(n89), .B1(n1), .Y(n94) );
  OAI31XL U52 ( .A0(n114), .A1(n2), .A2(n16), .B0(n90), .Y(n91) );
  OAI21XL U53 ( .A0(n81), .A1(n10), .B0(n5), .Y(n90) );
  NAND2X1 U54 ( .A(n8), .B(n2), .Y(n137) );
  OAI31XL U56 ( .A0(n101), .A1(n3), .A2(addr[2]), .B0(n113), .Y(n92) );
  OAI211X1 U58 ( .A0(n139), .A1(n83), .B0(n138), .C0(n137), .Y(n143) );
  NAND3X1 U59 ( .A(n82), .B(n83), .C(addr[6]), .Y(n138) );
  AOI2BB2X1 U65 ( .B0(n5), .B1(n16), .A0N(n6), .A1N(n136), .Y(n139) );
  OAI22XL U66 ( .A0(addr[5]), .A1(n133), .B0(n3), .B1(n132), .Y(n134) );
  OAI2BB2XL U68 ( .B0(n112), .B1(n122), .A0N(n1), .A1N(n99), .Y(n100) );
  OAI211X1 U69 ( .A0(n146), .A1(n2), .B0(n137), .C0(n113), .Y(n99) );
  NAND3X1 U70 ( .A(n5), .B(n82), .C(n3), .Y(n87) );
  AOI2BB2XL U71 ( .B0(n3), .B1(n105), .A0N(n137), .A1N(n132), .Y(n108) );
  OAI211XL U72 ( .A0(n104), .A1(n146), .B0(n103), .C0(n111), .Y(n105) );
  NAND3XL U73 ( .A(addr[5]), .B(n82), .C(n7), .Y(n103) );
  OAI22XL U74 ( .A0(n3), .A1(n114), .B0(n9), .B1(n115), .Y(n88) );
  NAND4X1 U75 ( .A(n110), .B(n109), .C(n108), .D(n107), .Y(dout[2]) );
  AOI32XL U76 ( .A0(addr[1]), .A1(addr[2]), .A2(n14), .B0(n100), .B1(n11), .Y(
        n110) );
  AOI221XL U77 ( .A0(n125), .A1(addr[4]), .B0(n141), .B1(n5), .C0(n106), .Y(
        n107) );
  AOI33XL U78 ( .A0(n5), .A1(n13), .A2(n2), .B0(n12), .B1(n146), .B2(n3), .Y(
        n145) );
  AOI222XL U79 ( .A0(n143), .A1(n11), .B0(n7), .B1(n142), .C0(n8), .C1(n141), 
        .Y(n144) );
  AOI32XL U80 ( .A0(n13), .A1(n6), .A2(n15), .B0(n4), .B1(n86), .Y(n97) );
  AOI22X1 U81 ( .A0(n7), .A1(n85), .B0(n2), .B1(n84), .Y(n98) );
  NAND2X1 U82 ( .A(n131), .B(n130), .Y(dout[3]) );
  AOI221XL U83 ( .A0(n120), .A1(n11), .B0(addr[2]), .B1(n119), .C0(n118), .Y(
        n131) );
  AOI211X1 U84 ( .A0(n13), .A1(n129), .B0(n128), .C0(n127), .Y(n130) );
  CLKINVX3 U85 ( .A(addr[2]), .Y(n11) );
  CLKINVX3 U86 ( .A(n3), .Y(n16) );
  CLKINVX3 U87 ( .A(n2), .Y(n82) );
endmodule


module sbox3_3 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134;

  NOR2X2 U35 ( .A(n7), .B(addr[3]), .Y(n109) );
  NOR2X2 U50 ( .A(addr[1]), .B(addr[6]), .Y(n108) );
  NOR2X2 U52 ( .A(n14), .B(n3), .Y(n88) );
  NOR2X2 U56 ( .A(n14), .B(n15), .Y(n95) );
  NOR2X1 U1 ( .A(n7), .B(n14), .Y(n107) );
  OAI221X1 U2 ( .A0(n125), .A1(n7), .B0(n4), .B1(addr[1]), .C0(n78), .Y(n105)
         );
  INVXL U3 ( .A(n2), .Y(n1) );
  NOR2X1 U4 ( .A(n20), .B(n4), .Y(n92) );
  NOR2X1 U5 ( .A(n9), .B(n4), .Y(n122) );
  NOR2X1 U6 ( .A(n78), .B(n4), .Y(n96) );
  CLKBUFX3 U7 ( .A(addr[2]), .Y(n4) );
  INVX1 U8 ( .A(addr[2]), .Y(n2) );
  NOR2X1 U9 ( .A(n4), .B(n3), .Y(n111) );
  BUFX4 U10 ( .A(addr[4]), .Y(n3) );
  OAI33X1 U11 ( .A0(n9), .A1(n126), .A2(n15), .B0(n7), .B1(n95), .B2(n120), 
        .Y(n80) );
  INVX3 U12 ( .A(n4), .Y(n15) );
  OAI221X1 U13 ( .A0(addr[5]), .A1(n91), .B0(n90), .B1(n17), .C0(n89), .Y(
        dout[1]) );
  NOR2X4 U14 ( .A(n76), .B(n79), .Y(n125) );
  NOR2X4 U15 ( .A(addr[3]), .B(n3), .Y(n131) );
  NOR2X4 U16 ( .A(n79), .B(addr[6]), .Y(n126) );
  INVX3 U17 ( .A(addr[1]), .Y(n79) );
  NAND2XL U18 ( .A(n95), .B(n125), .Y(n133) );
  OAI211XL U19 ( .A0(n3), .A1(n16), .B0(n129), .C0(n128), .Y(n130) );
  NAND4XL U20 ( .A(n115), .B(n114), .C(n113), .D(n112), .Y(n116) );
  CLKINVX1 U21 ( .A(n133), .Y(n13) );
  INVX1 U22 ( .A(n125), .Y(n18) );
  CLKINVX1 U23 ( .A(n107), .Y(n5) );
  NAND2X1 U24 ( .A(n20), .B(n6), .Y(n123) );
  CLKINVX1 U25 ( .A(n87), .Y(n6) );
  CLKINVX1 U26 ( .A(n121), .Y(n12) );
  CLKINVX1 U27 ( .A(n120), .Y(n19) );
  CLKINVX1 U28 ( .A(n115), .Y(n10) );
  CLKINVX1 U29 ( .A(n108), .Y(n78) );
  NOR2X1 U30 ( .A(n20), .B(n15), .Y(n104) );
  NOR2X1 U31 ( .A(n18), .B(n15), .Y(n110) );
  INVX1 U32 ( .A(n126), .Y(n77) );
  AOI21X1 U33 ( .A0(n14), .A1(n15), .B0(n95), .Y(n121) );
  OAI21XL U34 ( .A0(n111), .A1(n131), .B0(n125), .Y(n83) );
  CLKINVX1 U36 ( .A(n82), .Y(n20) );
  NOR2X1 U37 ( .A(n77), .B(n7), .Y(n87) );
  NOR2X1 U38 ( .A(n125), .B(n108), .Y(n120) );
  OAI21XL U39 ( .A0(n110), .A1(n92), .B0(n131), .Y(n101) );
  NAND2X1 U40 ( .A(n104), .B(n88), .Y(n115) );
  CLKINVX1 U41 ( .A(n88), .Y(n9) );
  CLKINVX1 U42 ( .A(n92), .Y(n16) );
  CLKINVX1 U43 ( .A(n111), .Y(n11) );
  CLKINVX1 U44 ( .A(n122), .Y(n8) );
  OR2X1 U45 ( .A(n104), .B(n96), .Y(n127) );
  OAI221X1 U46 ( .A0(n77), .A1(n11), .B0(n15), .B1(n6), .C0(n94), .Y(n99) );
  AOI221XL U47 ( .A0(n96), .A1(n3), .B0(n93), .B1(n7), .C0(n13), .Y(n94) );
  OAI21XL U48 ( .A0(n15), .A1(n78), .B0(n16), .Y(n93) );
  XNOR2X1 U49 ( .A(addr[5]), .B(addr[3]), .Y(n103) );
  CLKINVX1 U51 ( .A(addr[5]), .Y(n17) );
  OAI221X1 U53 ( .A0(n78), .A1(n11), .B0(n18), .B1(n9), .C0(n106), .Y(n117) );
  AOI221XL U54 ( .A0(addr[3]), .A1(n105), .B0(n104), .B1(n131), .C0(n13), .Y(
        n106) );
  CLKINVX1 U55 ( .A(addr[6]), .Y(n76) );
  NAND3X1 U57 ( .A(n4), .B(n79), .C(n109), .Y(n114) );
  NOR2X1 U58 ( .A(n76), .B(addr[1]), .Y(n82) );
  AOI32XL U59 ( .A0(n15), .A1(n14), .A2(n125), .B0(n124), .B1(n76), .Y(n129)
         );
  AOI22XL U60 ( .A0(n3), .A1(n127), .B0(n126), .B1(n131), .Y(n128) );
  OAI22XL U61 ( .A0(n3), .A1(n2), .B0(n4), .B1(n5), .Y(n124) );
  AOI222XL U62 ( .A0(n111), .A1(n126), .B0(n110), .B1(n14), .C0(n109), .C1(
        n108), .Y(n112) );
  OAI211XL U63 ( .A0(n107), .A1(n131), .B0(n2), .C0(addr[6]), .Y(n113) );
  OAI21XL U64 ( .A0(n1), .A1(addr[1]), .B0(n77), .Y(n81) );
  AOI221XL U65 ( .A0(n87), .A1(n14), .B0(n88), .B1(n126), .C0(n86), .Y(n90) );
  OAI211X1 U66 ( .A0(n85), .A1(n15), .B0(n84), .C0(n83), .Y(n86) );
  AOI222XL U67 ( .A0(n82), .A1(n14), .B0(n108), .B1(n107), .C0(n131), .C1(n79), 
        .Y(n85) );
  OAI21XL U68 ( .A0(n92), .A1(n13), .B0(addr[4]), .Y(n84) );
  AOI221XL U69 ( .A0(n126), .A1(n12), .B0(addr[3]), .B1(n127), .C0(n97), .Y(
        n98) );
  OAI22X1 U70 ( .A0(n18), .A1(n8), .B0(n5), .B1(n20), .Y(n97) );
  OAI211X1 U71 ( .A0(n78), .A1(n8), .B0(n119), .C0(n118), .Y(dout[3]) );
  AOI32XL U72 ( .A0(n126), .A1(n4), .A2(n103), .B0(n109), .B1(n110), .Y(n119)
         );
  AOI22XL U73 ( .A0(n117), .A1(n17), .B0(addr[5]), .B1(n116), .Y(n118) );
  AOI221XL U74 ( .A0(n122), .A1(n126), .B0(n96), .B1(n109), .C0(n10), .Y(n89)
         );
  AOI221XL U75 ( .A0(n131), .A1(n81), .B0(n95), .B1(n123), .C0(n80), .Y(n91)
         );
  NAND4X1 U76 ( .A(n102), .B(n114), .C(n101), .D(n100), .Y(dout[2]) );
  NAND3XL U77 ( .A(n3), .B(n125), .C(n103), .Y(n102) );
  AOI2BB2XL U78 ( .B0(addr[5]), .B1(n99), .A0N(addr[5]), .A1N(n98), .Y(n100)
         );
  OAI221X1 U79 ( .A0(n134), .A1(n17), .B0(n3), .B1(n133), .C0(n132), .Y(
        dout[4]) );
  AOI32XL U80 ( .A0(n131), .A1(n76), .A2(n1), .B0(n130), .B1(n17), .Y(n132) );
  AOI222XL U81 ( .A0(n12), .A1(n123), .B0(n122), .B1(addr[1]), .C0(n121), .C1(
        n19), .Y(n134) );
  CLKINVX3 U82 ( .A(n3), .Y(n7) );
  CLKINVX3 U83 ( .A(addr[3]), .Y(n14) );
endmodule


module sbox4_3 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126;

  OAI32X4 U12 ( .A0(n6), .A1(n2), .A2(addr[2]), .B0(n72), .B1(n108), .Y(n123)
         );
  OAI222X4 U20 ( .A0(addr[2]), .A1(n92), .B0(n106), .B1(n91), .C0(n90), .C1(
        n71), .Y(dout[2]) );
  OAI222X4 U33 ( .A0(addr[4]), .A1(n106), .B0(n16), .B1(n108), .C0(n2), .C1(
        n118), .Y(n83) );
  NAND2X2 U34 ( .A(addr[4]), .B(n2), .Y(n108) );
  NOR2X2 U43 ( .A(n8), .B(addr[4]), .Y(n113) );
  NOR2X2 U45 ( .A(n72), .B(n2), .Y(n111) );
  NAND2X2 U51 ( .A(n16), .B(n13), .Y(n118) );
  NOR2X2 U52 ( .A(n7), .B(addr[5]), .Y(n97) );
  NAND2X2 U53 ( .A(addr[6]), .B(addr[1]), .Y(n85) );
  NAND2X2 U54 ( .A(addr[1]), .B(n13), .Y(n116) );
  NOR2X2 U55 ( .A(n115), .B(n72), .Y(n121) );
  NAND2X2 U56 ( .A(n8), .B(n7), .Y(n115) );
  NAND2X2 U57 ( .A(addr[5]), .B(n7), .Y(n96) );
  NAND2X2 U58 ( .A(addr[6]), .B(n16), .Y(n106) );
  OAI222X1 U1 ( .A0(n6), .A1(n85), .B0(n97), .B1(n116), .C0(n7), .C1(n118), 
        .Y(n73) );
  CLKINVX1 U2 ( .A(n116), .Y(n12) );
  OAI31X4 U3 ( .A0(n118), .A1(n72), .A2(n7), .B0(n117), .Y(n119) );
  CLKINVX1 U4 ( .A(n8), .Y(n1) );
  CLKBUFX3 U5 ( .A(addr[3]), .Y(n2) );
  OAI221X1 U6 ( .A0(addr[2]), .A1(n80), .B0(n118), .B1(n105), .C0(n79), .Y(
        dout[1]) );
  INVX4 U7 ( .A(addr[5]), .Y(n72) );
  OAI31X1 U8 ( .A0(n108), .A1(addr[5]), .A2(n14), .B0(n107), .Y(n109) );
  AOI222XL U9 ( .A0(n7), .A1(n13), .B0(n113), .B1(n16), .C0(addr[1]), .C1(n8), 
        .Y(n114) );
  OAI222X1 U10 ( .A0(addr[1]), .A1(n84), .B0(n85), .B1(n74), .C0(n8), .C1(n107), .Y(n75) );
  NAND2XL U11 ( .A(n1), .B(addr[5]), .Y(n84) );
  AOI211XL U13 ( .A0(n83), .A1(n72), .B0(n82), .C0(n5), .Y(n92) );
  NAND2XL U14 ( .A(n7), .B(n72), .Y(n74) );
  CLKINVX1 U15 ( .A(n118), .Y(n10) );
  CLKINVX1 U16 ( .A(n115), .Y(n4) );
  CLKINVX1 U17 ( .A(n112), .Y(n11) );
  OAI21X1 U18 ( .A0(n12), .A1(n14), .B0(n71), .Y(n112) );
  AOI22X1 U19 ( .A0(n15), .A1(n111), .B0(n14), .B1(n113), .Y(n93) );
  OAI211X1 U21 ( .A0(n16), .A1(n115), .B0(n93), .C0(n3), .Y(n94) );
  CLKINVX1 U22 ( .A(n85), .Y(n15) );
  NAND2X1 U23 ( .A(n97), .B(n8), .Y(n105) );
  NAND2X1 U24 ( .A(n113), .B(n10), .Y(n98) );
  NAND2X1 U25 ( .A(n12), .B(n97), .Y(n107) );
  NAND2X1 U26 ( .A(n118), .B(n85), .Y(n110) );
  OAI21XL U27 ( .A0(n4), .A1(n72), .B0(n108), .Y(n95) );
  CLKINVX1 U28 ( .A(n84), .Y(n9) );
  CLKINVX1 U29 ( .A(addr[2]), .Y(n71) );
  OAI31X1 U30 ( .A0(n7), .A1(addr[6]), .A2(n72), .B0(n87), .Y(n88) );
  OAI21XL U31 ( .A0(n113), .A1(n6), .B0(n15), .Y(n87) );
  OAI211X1 U32 ( .A0(n76), .A1(n7), .B0(n98), .C0(n3), .Y(n77) );
  AOI222XL U35 ( .A0(addr[5]), .A1(addr[6]), .B0(n111), .B1(addr[1]), .C0(n14), 
        .C1(n2), .Y(n76) );
  NAND3XL U36 ( .A(n15), .B(n8), .C(addr[4]), .Y(n117) );
  OAI22XL U37 ( .A0(n116), .A1(n115), .B0(n1), .B1(n112), .Y(n78) );
  CLKINVX3 U38 ( .A(addr[4]), .Y(n7) );
  OAI2BB2XL U39 ( .B0(n115), .B1(n106), .A0N(n72), .A1N(n86), .Y(n89) );
  OAI221XL U40 ( .A0(n116), .A1(addr[4]), .B0(n108), .B1(addr[1]), .C0(n117), 
        .Y(n86) );
  CLKINVX1 U41 ( .A(addr[6]), .Y(n13) );
  CLKINVX1 U42 ( .A(n81), .Y(n5) );
  OAI21XL U44 ( .A0(n96), .A1(n118), .B0(n93), .Y(n82) );
  NAND3X1 U46 ( .A(n101), .B(n100), .C(n99), .Y(n102) );
  AOI32X1 U47 ( .A0(n96), .A1(n8), .A2(n12), .B0(n15), .B1(n95), .Y(n101) );
  AOI2BB2XL U48 ( .B0(n16), .B1(n121), .A0N(n98), .A1N(addr[5]), .Y(n99) );
  OAI21XL U49 ( .A0(n97), .A1(n6), .B0(n14), .Y(n100) );
  AOI2BB2XL U50 ( .B0(n14), .B1(n123), .A0N(n122), .A1N(n71), .Y(n124) );
  AOI211XL U59 ( .A0(n14), .A1(n121), .B0(n120), .C0(n119), .Y(n122) );
  OAI22XL U60 ( .A0(n116), .A1(n115), .B0(addr[5]), .B1(n114), .Y(n120) );
  CLKINVX1 U61 ( .A(n75), .Y(n3) );
  AOI32XL U62 ( .A0(n12), .A1(n96), .A2(n1), .B0(addr[1]), .B1(n121), .Y(n81)
         );
  AOI222XL U63 ( .A0(n14), .A1(n6), .B0(n121), .B1(n116), .C0(n2), .C1(n73), 
        .Y(n80) );
  AOI22XL U64 ( .A0(n78), .A1(n72), .B0(addr[2]), .B1(n77), .Y(n79) );
  NAND2XL U65 ( .A(n111), .B(addr[4]), .Y(n91) );
  AOI211X1 U66 ( .A0(n9), .A1(n110), .B0(n89), .C0(n88), .Y(n90) );
  OAI211X1 U67 ( .A0(n106), .A1(n105), .B0(n104), .C0(n103), .Y(dout[3]) );
  AOI32X1 U68 ( .A0(n2), .A1(n6), .A2(n12), .B0(n94), .B1(n71), .Y(n104) );
  AOI22XL U69 ( .A0(addr[2]), .A1(n102), .B0(n10), .B1(n123), .Y(n103) );
  OAI211X1 U70 ( .A0(addr[2]), .A1(n126), .B0(n125), .C0(n124), .Y(dout[4]) );
  AOI32X1 U71 ( .A0(n15), .A1(n6), .A2(n2), .B0(n11), .B1(n9), .Y(n125) );
  AOI221XL U72 ( .A0(n10), .A1(n111), .B0(n4), .B1(n110), .C0(n109), .Y(n126)
         );
  CLKINVX3 U73 ( .A(n96), .Y(n6) );
  CLKINVX3 U74 ( .A(n2), .Y(n8) );
  CLKINVX3 U75 ( .A(n106), .Y(n14) );
  CLKINVX3 U76 ( .A(addr[1]), .Y(n16) );
endmodule


module sbox5_3 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121;

  OAI222X4 U18 ( .A0(addr[3]), .A1(n106), .B0(n14), .B1(n90), .C0(n5), .C1(n70), .Y(n93) );
  OAI22X2 U40 ( .A0(addr[5]), .A1(n106), .B0(n68), .B1(n114), .Y(n116) );
  NOR2X2 U41 ( .A(n3), .B(addr[3]), .Y(n102) );
  NAND2X2 U45 ( .A(addr[6]), .B(n70), .Y(n114) );
  NAND2X2 U50 ( .A(n70), .B(n14), .Y(n110) );
  NAND2X2 U52 ( .A(addr[1]), .B(n14), .Y(n113) );
  NAND2X2 U54 ( .A(addr[1]), .B(addr[6]), .Y(n106) );
  NAND2X2 U55 ( .A(addr[3]), .B(n5), .Y(n121) );
  OAI221X4 U1 ( .A0(n111), .A1(n110), .B0(n121), .B1(n114), .C0(n109), .Y(n112) );
  OAI221X4 U2 ( .A0(n107), .A1(n121), .B0(n111), .B1(n113), .C0(n85), .Y(n86)
         );
  OAI31X1 U3 ( .A0(n9), .A1(addr[5]), .A2(addr[1]), .B0(n81), .Y(n73) );
  CLKINVX1 U4 ( .A(addr[5]), .Y(n1) );
  OAI221X4 U5 ( .A0(n5), .A1(n114), .B0(n68), .B1(n113), .C0(n120), .Y(n115)
         );
  AOI221XL U6 ( .A0(n93), .A1(n1), .B0(n15), .B1(n7), .C0(n92), .Y(n105) );
  INVX3 U7 ( .A(addr[5]), .Y(n68) );
  OAI32X1 U8 ( .A0(n114), .A1(addr[5]), .A2(n3), .B0(n4), .B1(n107), .Y(n79)
         );
  AOI32XL U9 ( .A0(n7), .A1(n98), .A2(n13), .B0(n2), .B1(n73), .Y(n77) );
  CLKBUFX3 U10 ( .A(addr[4]), .Y(n2) );
  CLKINVX1 U11 ( .A(n81), .Y(n6) );
  NAND2X1 U12 ( .A(n16), .B(n7), .Y(n81) );
  CLKINVX1 U13 ( .A(n110), .Y(n11) );
  CLKXOR2X2 U14 ( .A(n9), .B(n68), .Y(n94) );
  AOI2BB1X1 U15 ( .A0N(n5), .A1N(n1), .B0(n7), .Y(n111) );
  NOR2X1 U16 ( .A(n121), .B(n68), .Y(n91) );
  NOR2BX1 U17 ( .AN(n116), .B(n90), .Y(n83) );
  NAND2X1 U19 ( .A(n11), .B(n68), .Y(n120) );
  CLKINVX1 U20 ( .A(n113), .Y(n13) );
  NAND2X1 U21 ( .A(n13), .B(n68), .Y(n107) );
  CLKINVX1 U22 ( .A(n121), .Y(n4) );
  OAI31X1 U23 ( .A0(n69), .A1(n7), .A2(n113), .B0(n99), .Y(n72) );
  CLKINVX1 U24 ( .A(n106), .Y(n15) );
  OAI2BB2XL U25 ( .B0(n1), .B1(n113), .A0N(n98), .A1N(n16), .Y(n101) );
  CLKINVX1 U26 ( .A(n114), .Y(n16) );
  CLKINVX1 U27 ( .A(n90), .Y(n8) );
  CLKINVX1 U28 ( .A(addr[1]), .Y(n70) );
  CLKINVX1 U29 ( .A(addr[3]), .Y(n9) );
  CLKINVX1 U30 ( .A(addr[6]), .Y(n14) );
  AOI211X1 U31 ( .A0(n91), .A1(addr[1]), .B0(n80), .C0(n79), .Y(n89) );
  OAI2BB2XL U32 ( .B0(n111), .B1(n106), .A0N(n94), .A1N(n11), .Y(n80) );
  AOI211X1 U33 ( .A0(n102), .A1(n84), .B0(n83), .C0(n82), .Y(n85) );
  OAI21XL U34 ( .A0(n14), .A1(n1), .B0(n106), .Y(n84) );
  NOR3XL U35 ( .A(n94), .B(n3), .C(n110), .Y(n82) );
  AOI222XL U36 ( .A0(n15), .A1(n8), .B0(addr[5]), .B1(n108), .C0(n12), .C1(n5), 
        .Y(n109) );
  CLKINVX1 U37 ( .A(n107), .Y(n12) );
  OAI21XL U38 ( .A0(addr[6]), .A1(addr[3]), .B0(n106), .Y(n108) );
  NAND2X1 U39 ( .A(addr[3]), .B(n3), .Y(n90) );
  NAND2X1 U42 ( .A(n2), .B(addr[5]), .Y(n98) );
  NAND2X1 U43 ( .A(n3), .B(n9), .Y(n97) );
  OAI21XL U44 ( .A0(addr[1]), .A1(n97), .B0(n96), .Y(n103) );
  AOI33XL U46 ( .A0(n3), .A1(n95), .A2(addr[5]), .B0(n94), .B1(n5), .B2(
        addr[1]), .Y(n96) );
  OAI21XL U47 ( .A0(n70), .A1(n9), .B0(n114), .Y(n95) );
  OAI21XL U48 ( .A0(addr[6]), .A1(n121), .B0(n99), .Y(n100) );
  NAND2X1 U49 ( .A(n71), .B(n11), .Y(n99) );
  XOR2X1 U51 ( .A(n69), .B(n3), .Y(n71) );
  AOI2BB2XL U53 ( .B0(n102), .B1(n116), .A0N(n2), .A1N(n75), .Y(n76) );
  AOI211X1 U56 ( .A0(n10), .A1(n3), .B0(n74), .C0(n83), .Y(n75) );
  AO22XL U57 ( .A0(n13), .A1(n4), .B0(addr[6]), .B1(n102), .Y(n74) );
  CLKINVX1 U58 ( .A(n120), .Y(n10) );
  CLKINVX1 U59 ( .A(n2), .Y(n69) );
  AO22XL U60 ( .A0(n13), .A1(n8), .B0(addr[6]), .B1(n91), .Y(n92) );
  AOI222XL U61 ( .A0(n116), .A1(n5), .B0(addr[3]), .B1(n115), .C0(n13), .C1(n7), .Y(n117) );
  OAI221X1 U62 ( .A0(n2), .A1(n105), .B0(n110), .B1(n121), .C0(n104), .Y(
        dout[3]) );
  AOI222XL U63 ( .A0(n2), .A1(n103), .B0(n102), .B1(n101), .C0(n100), .C1(n1), 
        .Y(n104) );
  OAI211X1 U64 ( .A0(n2), .A1(n89), .B0(n88), .C0(n87), .Y(dout[2]) );
  AOI33XL U65 ( .A0(n4), .A1(n98), .A2(n16), .B0(n3), .B1(n94), .B2(n11), .Y(
        n88) );
  AOI222XL U66 ( .A0(n6), .A1(n68), .B0(n2), .B1(n86), .C0(n91), .C1(n15), .Y(
        n87) );
  OAI211X1 U67 ( .A0(n78), .A1(n68), .B0(n77), .C0(n76), .Y(dout[1]) );
  AOI221XL U68 ( .A0(n4), .A1(addr[1]), .B0(n15), .B1(n7), .C0(n72), .Y(n78)
         );
  OAI211X1 U69 ( .A0(n121), .A1(n120), .B0(n119), .C0(n118), .Y(dout[4]) );
  AOI32XL U70 ( .A0(n7), .A1(n114), .A2(addr[5]), .B0(n2), .B1(n112), .Y(n119)
         );
  AOI2BB2X1 U71 ( .B0(n6), .B1(n68), .A0N(n2), .A1N(n117), .Y(n118) );
  BUFX4 U72 ( .A(addr[2]), .Y(n3) );
  CLKINVX3 U73 ( .A(n3), .Y(n5) );
  CLKINVX3 U74 ( .A(n97), .Y(n7) );
endmodule


module sbox6_3 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147;

  NAND2X2 U39 ( .A(n138), .B(addr[3]), .Y(n147) );
  NOR2X2 U47 ( .A(n15), .B(n13), .Y(n138) );
  NOR2X2 U50 ( .A(n81), .B(n4), .Y(n119) );
  NOR2X2 U58 ( .A(n84), .B(n81), .Y(n125) );
  NAND2X2 U61 ( .A(n97), .B(n103), .Y(n112) );
  NOR2X2 U62 ( .A(n11), .B(addr[1]), .Y(n103) );
  NOR2X2 U63 ( .A(n84), .B(addr[3]), .Y(n97) );
  NAND2X2 U64 ( .A(n117), .B(n131), .Y(n140) );
  NOR2X2 U65 ( .A(n5), .B(addr[3]), .Y(n131) );
  NOR2X2 U66 ( .A(n83), .B(addr[6]), .Y(n117) );
  NOR2X1 U1 ( .A(n15), .B(addr[3]), .Y(n102) );
  OAI222X1 U2 ( .A0(n91), .A1(n85), .B0(n3), .B1(n82), .C0(addr[5]), .C1(n17), 
        .Y(n92) );
  CLKINVX1 U3 ( .A(n84), .Y(n1) );
  INVX4 U4 ( .A(n4), .Y(n84) );
  CLKBUFX3 U5 ( .A(addr[4]), .Y(n4) );
  CLKINVX1 U6 ( .A(addr[3]), .Y(n2) );
  INVX3 U7 ( .A(addr[3]), .Y(n81) );
  OAI221X1 U8 ( .A0(n11), .A1(n18), .B0(n81), .B1(n8), .C0(n86), .Y(n90) );
  INVX2 U9 ( .A(n96), .Y(n8) );
  CLKINVX1 U10 ( .A(n15), .Y(n3) );
  BUFX4 U11 ( .A(addr[2]), .Y(n5) );
  NOR2X4 U12 ( .A(addr[1]), .B(addr[6]), .Y(n130) );
  OAI22X1 U13 ( .A0(n81), .A1(n11), .B0(addr[1]), .B1(n17), .Y(n142) );
  OAI221X4 U14 ( .A0(n123), .A1(n10), .B0(n13), .B1(n85), .C0(n7), .Y(n124) );
  NOR2X4 U15 ( .A(n5), .B(addr[5]), .Y(n143) );
  INVX1 U16 ( .A(n130), .Y(n14) );
  CLKINVX1 U17 ( .A(n125), .Y(n18) );
  NAND2X1 U18 ( .A(n14), .B(n8), .Y(n105) );
  INVXL U19 ( .A(n121), .Y(n16) );
  CLKINVX1 U20 ( .A(n138), .Y(n12) );
  AOI211X1 U21 ( .A0(n85), .A1(n81), .B0(n131), .C0(n143), .Y(n121) );
  CLKINVX1 U22 ( .A(n117), .Y(n13) );
  CLKINVX1 U23 ( .A(n119), .Y(n17) );
  NOR2X1 U24 ( .A(n8), .B(n123), .Y(n144) );
  NOR2X1 U25 ( .A(n83), .B(n11), .Y(n96) );
  CLKINVX1 U26 ( .A(n103), .Y(n10) );
  OAI211X1 U27 ( .A0(n14), .A1(n18), .B0(n104), .C0(n112), .Y(n108) );
  OAI21XL U28 ( .A0(n103), .A1(n117), .B0(n102), .Y(n104) );
  OAI21XL U29 ( .A0(n132), .A1(n11), .B0(n2), .Y(n86) );
  AOI21X1 U30 ( .A0(n84), .A1(n102), .B0(n125), .Y(n91) );
  OAI2BB2XL U31 ( .B0(n143), .B1(n14), .A0N(n143), .A1N(n117), .Y(n118) );
  CLKINVX1 U32 ( .A(n122), .Y(n7) );
  CLKINVX1 U33 ( .A(n126), .Y(n9) );
  CLKINVX1 U34 ( .A(n97), .Y(n82) );
  NAND2BX1 U35 ( .AN(n144), .B(n137), .Y(n107) );
  CLKINVX1 U36 ( .A(addr[1]), .Y(n83) );
  NOR2X1 U37 ( .A(n8), .B(n3), .Y(n122) );
  NOR2X1 U38 ( .A(addr[1]), .B(n1), .Y(n132) );
  OAI22X1 U40 ( .A0(n17), .A1(n13), .B0(n5), .B1(n9), .Y(n88) );
  NAND2X1 U41 ( .A(n5), .B(n85), .Y(n123) );
  NAND4X1 U42 ( .A(n147), .B(n140), .C(n100), .D(n99), .Y(n101) );
  AOI222XL U43 ( .A0(n98), .A1(n15), .B0(n102), .B1(n130), .C0(n97), .C1(n105), 
        .Y(n99) );
  NAND3X1 U44 ( .A(n5), .B(n17), .C(n96), .Y(n100) );
  OAI221X1 U45 ( .A0(n81), .A1(n10), .B0(n17), .B1(n11), .C0(n9), .Y(n98) );
  AOI22X1 U46 ( .A0(n4), .A1(n115), .B0(addr[5]), .B1(n114), .Y(n129) );
  OAI21XL U48 ( .A0(n121), .A1(n14), .B0(n147), .Y(n115) );
  OAI21XL U49 ( .A0(n113), .A1(n15), .B0(n112), .Y(n114) );
  AOI221XL U51 ( .A0(n119), .A1(n83), .B0(n130), .B1(addr[3]), .C0(n111), .Y(
        n113) );
  OAI22XL U52 ( .A0(n13), .A1(n84), .B0(addr[3]), .B1(n8), .Y(n111) );
  AOI211X1 U53 ( .A0(n4), .A1(n135), .B0(n134), .C0(n133), .Y(n136) );
  OA21XL U54 ( .A0(n2), .A1(n3), .B0(n132), .Y(n133) );
  OAI2BB2XL U55 ( .B0(n1), .B1(n7), .A0N(n131), .A1N(n130), .Y(n134) );
  OAI22X1 U56 ( .A0(n5), .A1(n13), .B0(n15), .B1(n8), .Y(n135) );
  CLKINVX3 U57 ( .A(addr[5]), .Y(n85) );
  AOI2BB2X1 U59 ( .B0(n5), .B1(n130), .A0N(n3), .A1N(n10), .Y(n137) );
  NOR2X1 U60 ( .A(n10), .B(n1), .Y(n126) );
  AOI2BB2XL U67 ( .B0(n143), .B1(n90), .A0N(n89), .A1N(n85), .Y(n94) );
  AOI211X1 U68 ( .A0(n122), .A1(n4), .B0(n88), .C0(n87), .Y(n89) );
  OAI32X1 U69 ( .A0(n10), .A1(n81), .A2(n15), .B0(n12), .B1(n82), .Y(n87) );
  NAND3X1 U70 ( .A(n147), .B(n140), .C(n139), .Y(n141) );
  AOI32X1 U71 ( .A0(n5), .A1(n83), .A2(n4), .B0(n138), .B1(n84), .Y(n139) );
  AO22XL U72 ( .A0(n143), .A1(n1), .B0(n116), .B1(n84), .Y(n120) );
  OAI21XL U73 ( .A0(n3), .A1(n85), .B0(n123), .Y(n116) );
  CLKINVX1 U74 ( .A(n106), .Y(n6) );
  AOI32XL U75 ( .A0(n105), .A1(n84), .A2(n2), .B0(addr[1]), .B1(n125), .Y(n106) );
  OAI211X1 U76 ( .A0(n84), .A1(n140), .B0(n110), .C0(n109), .Y(dout[2]) );
  AOI222XL U77 ( .A0(n108), .A1(n85), .B0(n143), .B1(n6), .C0(n119), .C1(n107), 
        .Y(n109) );
  AOI2BB2XL U78 ( .B0(addr[5]), .B1(n101), .A0N(n15), .A1N(n112), .Y(n110) );
  OAI211X1 U79 ( .A0(n1), .A1(n147), .B0(n146), .C0(n145), .Y(dout[4]) );
  AOI222XL U80 ( .A0(n144), .A1(n81), .B0(n143), .B1(n142), .C0(n141), .C1(n85), .Y(n145) );
  OA22X1 U81 ( .A0(n18), .A1(n137), .B0(n136), .B1(n85), .Y(n146) );
  NAND3X1 U82 ( .A(n129), .B(n128), .C(n127), .Y(dout[3]) );
  AOI32XL U83 ( .A0(n120), .A1(n81), .A2(addr[1]), .B0(n119), .B1(n118), .Y(
        n128) );
  AOI222XL U84 ( .A0(n144), .A1(n84), .B0(n126), .B1(n16), .C0(n125), .C1(n124), .Y(n127) );
  NAND3BX1 U85 ( .AN(n95), .B(n94), .C(n93), .Y(dout[1]) );
  OAI222X1 U86 ( .A0(n140), .A1(n4), .B0(n112), .B1(n15), .C0(n8), .C1(n91), 
        .Y(n95) );
  AOI32XL U87 ( .A0(addr[1]), .A1(n85), .A2(n125), .B0(n130), .B1(n92), .Y(n93) );
  CLKINVX3 U88 ( .A(addr[6]), .Y(n11) );
  CLKINVX3 U89 ( .A(n5), .Y(n15) );
endmodule


module sbox7_3 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148;

  OAI222X4 U19 ( .A0(n20), .A1(n129), .B0(n4), .B1(n13), .C0(addr[1]), .C1(n12), .Y(n122) );
  OAI33X4 U33 ( .A0(addr[1]), .A1(n4), .A2(n5), .B0(n18), .B1(n21), .B2(n6), 
        .Y(n97) );
  NOR2X2 U44 ( .A(n10), .B(n4), .Y(n116) );
  NOR2X2 U48 ( .A(addr[1]), .B(addr[6]), .Y(n136) );
  NOR2X2 U51 ( .A(n87), .B(n10), .Y(n125) );
  NOR2X2 U52 ( .A(n18), .B(addr[3]), .Y(n131) );
  NOR2X2 U58 ( .A(n93), .B(n124), .Y(n142) );
  NOR2X2 U60 ( .A(n19), .B(addr[1]), .Y(n93) );
  NOR2X2 U62 ( .A(n84), .B(n3), .Y(n137) );
  NOR2X2 U65 ( .A(n19), .B(n86), .Y(n140) );
  NAND2X1 U1 ( .A(n3), .B(n4), .Y(n119) );
  CLKBUFX3 U2 ( .A(addr[4]), .Y(n4) );
  CLKINVX1 U3 ( .A(n84), .Y(n1) );
  CLKINVX1 U4 ( .A(n21), .Y(n2) );
  CLKBUFX3 U5 ( .A(addr[2]), .Y(n5) );
  OAI31X1 U6 ( .A0(n10), .A1(n84), .A2(n86), .B0(n117), .Y(n121) );
  NOR2X4 U7 ( .A(n86), .B(addr[6]), .Y(n124) );
  OAI22X1 U8 ( .A0(addr[1]), .A1(n12), .B0(n5), .B1(n113), .Y(n100) );
  OAI22X1 U9 ( .A0(n4), .A1(n87), .B0(addr[3]), .B1(n83), .Y(n103) );
  AOI211XL U10 ( .A0(n5), .A1(n17), .B0(n131), .C0(n130), .Y(n132) );
  NOR3XL U11 ( .A(n20), .B(addr[3]), .C(n2), .Y(n130) );
  OAI21XL U12 ( .A0(n3), .A1(n1), .B0(n119), .Y(n89) );
  BUFX4 U13 ( .A(addr[5]), .Y(n3) );
  AOI221XL U14 ( .A0(n140), .A1(n89), .B0(n109), .B1(n17), .C0(n88), .Y(n96)
         );
  CLKINVX1 U15 ( .A(n140), .Y(n18) );
  OAI2BB2XL U16 ( .B0(n142), .B1(n83), .A0N(n141), .A1N(n140), .Y(n143) );
  CLKINVX1 U17 ( .A(n125), .Y(n8) );
  CLKINVX1 U18 ( .A(n142), .Y(n17) );
  NAND2X1 U20 ( .A(n8), .B(n14), .Y(n105) );
  CLKINVX1 U21 ( .A(n123), .Y(n11) );
  CLKINVX1 U22 ( .A(n109), .Y(n9) );
  NAND2X1 U23 ( .A(n124), .B(n10), .Y(n113) );
  CLKINVX1 U24 ( .A(n137), .Y(n83) );
  NOR2X1 U25 ( .A(n83), .B(n10), .Y(n109) );
  CLKINVX1 U26 ( .A(n136), .Y(n20) );
  OAI22XL U27 ( .A0(n137), .A1(n13), .B0(n86), .B1(n9), .Y(n146) );
  OAI21X1 U28 ( .A0(n84), .A1(n8), .B0(n129), .Y(n141) );
  NAND2X1 U29 ( .A(n116), .B(n87), .Y(n129) );
  CLKINVX1 U30 ( .A(n93), .Y(n16) );
  OAI21XL U31 ( .A0(n119), .A1(n16), .B0(n118), .Y(n120) );
  OAI21XL U32 ( .A0(n125), .A1(n137), .B0(n124), .Y(n118) );
  NOR2X1 U34 ( .A(n87), .B(n12), .Y(n123) );
  CLKINVX1 U35 ( .A(n145), .Y(n12) );
  OAI22XL U36 ( .A0(n137), .A1(n113), .B0(n19), .B1(n11), .Y(n88) );
  CLKINVX1 U37 ( .A(n116), .Y(n6) );
  CLKINVX1 U38 ( .A(n131), .Y(n13) );
  CLKINVX1 U39 ( .A(n134), .Y(n14) );
  NOR2XL U40 ( .A(n125), .B(n84), .Y(n110) );
  CLKINVX1 U41 ( .A(n119), .Y(n85) );
  CLKINVX1 U42 ( .A(n103), .Y(n15) );
  OA21XL U43 ( .A0(n7), .A1(n16), .B0(n117), .Y(n102) );
  CLKINVX1 U45 ( .A(n105), .Y(n7) );
  OAI2BB1XL U46 ( .A0N(n103), .A1N(n124), .B0(n102), .Y(n104) );
  OAI22X1 U47 ( .A0(n87), .A1(n6), .B0(n4), .B1(n14), .Y(n112) );
  NOR4X1 U49 ( .A(n4), .B(addr[3]), .C(n86), .D(n21), .Y(n99) );
  XNOR2X1 U50 ( .A(addr[6]), .B(n5), .Y(n101) );
  AOI211X1 U53 ( .A0(n116), .A1(addr[6]), .B0(n115), .C0(n114), .Y(n128) );
  OAI222X1 U54 ( .A0(n111), .A1(n18), .B0(n110), .B1(n16), .C0(n20), .C1(n9), 
        .Y(n115) );
  OAI2BB2XL U55 ( .B0(n85), .B1(n113), .A0N(n86), .A1N(n112), .Y(n114) );
  OA21XL U56 ( .A0(n10), .A1(n3), .B0(n11), .Y(n111) );
  NAND2X1 U57 ( .A(n5), .B(n136), .Y(n133) );
  CLKINVX1 U59 ( .A(addr[6]), .Y(n19) );
  AOI211X1 U61 ( .A0(n131), .A1(n3), .B0(n92), .C0(n91), .Y(n95) );
  OAI221X1 U63 ( .A0(n86), .A1(n12), .B0(n18), .B1(n83), .C0(n102), .Y(n92) );
  OAI31X1 U64 ( .A0(n10), .A1(n84), .A2(n20), .B0(n90), .Y(n91) );
  AO21XL U66 ( .A0(n119), .A1(n129), .B0(addr[6]), .Y(n90) );
  NOR2X1 U67 ( .A(n84), .B(addr[3]), .Y(n145) );
  AOI21XL U68 ( .A0(addr[3]), .A1(n98), .B0(n97), .Y(n108) );
  OAI2BB1XL U69 ( .A0N(n21), .A1N(n124), .B0(n133), .Y(n98) );
  NAND3X1 U70 ( .A(n136), .B(n10), .C(n3), .Y(n117) );
  NOR2X1 U71 ( .A(addr[3]), .B(n3), .Y(n134) );
  OAI21X1 U72 ( .A0(n5), .A1(n142), .B0(n133), .Y(n138) );
  OAI22XL U73 ( .A0(n142), .A1(n6), .B0(n1), .B1(n132), .Y(n135) );
  AO21X1 U74 ( .A0(n139), .A1(n87), .B0(n138), .Y(n144) );
  OAI21XL U75 ( .A0(n2), .A1(n86), .B0(n16), .Y(n139) );
  OAI221X1 U76 ( .A0(n96), .A1(n21), .B0(n5), .B1(n95), .C0(n94), .Y(dout[1])
         );
  AOI2BB2X1 U77 ( .B0(n93), .B1(n112), .A0N(n133), .A1N(n15), .Y(n94) );
  OAI211X1 U78 ( .A0(n128), .A1(n21), .B0(n127), .C0(n126), .Y(dout[3]) );
  AOI32XL U79 ( .A0(n125), .A1(n1), .A2(n124), .B0(n123), .B1(n136), .Y(n126)
         );
  OAI31X1 U80 ( .A0(n122), .A1(n121), .A2(n120), .B0(n21), .Y(n127) );
  OAI221X1 U81 ( .A0(n3), .A1(n108), .B0(n107), .B1(n87), .C0(n106), .Y(
        dout[2]) );
  AOI32XL U82 ( .A0(n105), .A1(n21), .A2(n140), .B0(n2), .B1(n104), .Y(n106)
         );
  AOI211X1 U83 ( .A0(n101), .A1(n4), .B0(n100), .C0(n99), .Y(n107) );
  NAND2X1 U84 ( .A(n148), .B(n147), .Y(dout[4]) );
  AOI222XL U85 ( .A0(n136), .A1(n141), .B0(n3), .B1(n135), .C0(n134), .C1(n138), .Y(n148) );
  AOI222XL U86 ( .A0(n5), .A1(n146), .B0(n145), .B1(n144), .C0(n143), .C1(n21), 
        .Y(n147) );
  CLKINVX3 U87 ( .A(addr[3]), .Y(n10) );
  CLKINVX3 U88 ( .A(n5), .Y(n21) );
  CLKINVX3 U89 ( .A(n4), .Y(n84) );
  CLKINVX3 U90 ( .A(addr[1]), .Y(n86) );
  CLKINVX3 U91 ( .A(n3), .Y(n87) );
endmodule


module sbox8_3 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132;

  NAND2X2 U41 ( .A(addr[6]), .B(n10), .Y(n131) );
  NAND2X2 U48 ( .A(addr[4]), .B(n13), .Y(n123) );
  NAND2X2 U49 ( .A(n2), .B(n74), .Y(n87) );
  NAND2X2 U50 ( .A(addr[1]), .B(n6), .Y(n124) );
  NAND2X2 U54 ( .A(addr[2]), .B(n15), .Y(n116) );
  NAND2X2 U60 ( .A(addr[6]), .B(addr[1]), .Y(n105) );
  NAND2X2 U61 ( .A(n10), .B(n6), .Y(n108) );
  OAI32X1 U1 ( .A0(n6), .A1(addr[4]), .A2(n92), .B0(n115), .B1(n108), .Y(n96)
         );
  OAI31X1 U2 ( .A0(n123), .A1(addr[6]), .A2(n116), .B0(n109), .Y(n110) );
  AOI222X1 U3 ( .A0(n88), .A1(addr[2]), .B0(n74), .B1(n16), .C0(n75), .C1(n92), 
        .Y(n114) );
  OAI222X1 U4 ( .A0(addr[2]), .A1(n126), .B0(n13), .B1(n125), .C0(n124), .C1(
        n123), .Y(n127) );
  OAI221X1 U5 ( .A0(n105), .A1(n87), .B0(addr[4]), .B1(n108), .C0(n86), .Y(n90) );
  NAND2X4 U6 ( .A(addr[4]), .B(n2), .Y(n115) );
  AOI32XL U7 ( .A0(n4), .A1(n14), .A2(n2), .B0(n5), .B1(n117), .Y(n130) );
  OA21XL U8 ( .A0(n75), .A1(n15), .B0(n121), .Y(n78) );
  INVXL U9 ( .A(n119), .Y(n3) );
  INVX3 U10 ( .A(n2), .Y(n13) );
  BUFX4 U11 ( .A(addr[3]), .Y(n2) );
  CLKBUFX3 U12 ( .A(addr[5]), .Y(n1) );
  CLKINVX1 U13 ( .A(n108), .Y(n5) );
  CLKINVX1 U14 ( .A(n107), .Y(n11) );
  CLKINVX1 U15 ( .A(n93), .Y(n12) );
  NAND2X1 U16 ( .A(n13), .B(n74), .Y(n93) );
  NAND2X1 U17 ( .A(n75), .B(n15), .Y(n121) );
  OAI21XL U18 ( .A0(n115), .A1(n15), .B0(n107), .Y(n77) );
  OAI21X1 U19 ( .A0(n74), .A1(n15), .B0(n123), .Y(n88) );
  OAI31XL U20 ( .A0(n115), .A1(n10), .A2(n116), .B0(n118), .Y(n94) );
  CLKINVX1 U21 ( .A(n131), .Y(n9) );
  NAND2X1 U22 ( .A(n14), .B(n13), .Y(n107) );
  OAI22XL U23 ( .A0(n116), .A1(n123), .B0(n14), .B1(n115), .Y(n117) );
  OAI22XL U24 ( .A0(n123), .A1(n108), .B0(n131), .B1(n93), .Y(n95) );
  OAI2BB2XL U25 ( .B0(n115), .B1(n131), .A0N(n88), .A1N(n8), .Y(n89) );
  AOI211XL U26 ( .A0(n108), .A1(n105), .B0(n74), .C0(n121), .Y(n85) );
  CLKINVX1 U27 ( .A(n124), .Y(n4) );
  OAI22XL U28 ( .A0(n14), .A1(n123), .B0(n78), .B1(n87), .Y(n81) );
  NAND2BX2 U29 ( .AN(n78), .B(n13), .Y(n120) );
  NAND2XL U30 ( .A(n115), .B(n93), .Y(n104) );
  OAI2BB2XL U31 ( .B0(n106), .B1(n105), .A0N(n104), .A1N(n4), .Y(n111) );
  NOR2BXL U32 ( .AN(n123), .B(n103), .Y(n106) );
  NAND3X1 U33 ( .A(n104), .B(n10), .C(n14), .Y(n84) );
  AO21X1 U34 ( .A0(n14), .A1(n8), .B0(n101), .Y(n102) );
  OAI33X1 U35 ( .A0(n6), .A1(n13), .A2(n100), .B0(n75), .B1(n103), .B2(n124), 
        .Y(n101) );
  OA22XL U36 ( .A0(n107), .A1(n131), .B0(n120), .B1(n124), .Y(n98) );
  CLKINVX1 U37 ( .A(n125), .Y(n7) );
  OAI21XL U38 ( .A0(n4), .A1(n9), .B0(addr[4]), .Y(n86) );
  NAND2X1 U39 ( .A(n1), .B(n75), .Y(n100) );
  OAI221X1 U40 ( .A0(n124), .A1(n121), .B0(addr[1]), .B1(n120), .C0(n3), .Y(
        n128) );
  OAI31XL U42 ( .A0(n75), .A1(n10), .A2(n13), .B0(n118), .Y(n119) );
  NAND2X1 U43 ( .A(n8), .B(addr[2]), .Y(n125) );
  NAND4XL U44 ( .A(n9), .B(n1), .C(n2), .D(addr[2]), .Y(n109) );
  NAND3X1 U45 ( .A(n14), .B(n6), .C(n2), .Y(n118) );
  OAI21XL U46 ( .A0(n1), .A1(n87), .B0(n114), .Y(n76) );
  OAI22XL U47 ( .A0(n108), .A1(n120), .B0(n79), .B1(n100), .Y(n80) );
  AOI221XL U51 ( .A0(n9), .A1(n13), .B0(n8), .B1(n2), .C0(n91), .Y(n79) );
  NOR2X1 U52 ( .A(n1), .B(n2), .Y(n103) );
  NOR2X1 U53 ( .A(n87), .B(addr[6]), .Y(n91) );
  NOR2X1 U55 ( .A(n13), .B(n1), .Y(n92) );
  CLKINVX1 U56 ( .A(n100), .Y(n16) );
  OA21XL U57 ( .A0(n1), .A1(n115), .B0(n120), .Y(n132) );
  AOI221XL U58 ( .A0(n5), .A1(n2), .B0(n8), .B1(addr[4]), .C0(n122), .Y(n126)
         );
  OAI22XL U59 ( .A0(n2), .A1(n10), .B0(addr[4]), .B1(n131), .Y(n122) );
  OAI211X1 U62 ( .A0(addr[2]), .A1(n99), .B0(n98), .C0(n97), .Y(dout[2]) );
  AOI221XL U63 ( .A0(addr[2]), .A1(n96), .B0(n1), .B1(n95), .C0(n94), .Y(n97)
         );
  AOI221XL U64 ( .A0(n91), .A1(n1), .B0(n90), .B1(n15), .C0(n89), .Y(n99) );
  OAI211X1 U65 ( .A0(n132), .A1(n131), .B0(n130), .C0(n129), .Y(dout[4]) );
  AOI222XL U66 ( .A0(n128), .A1(n74), .B0(n1), .B1(n127), .C0(n11), .C1(n8), 
        .Y(n129) );
  OAI211X1 U67 ( .A0(addr[1]), .A1(n114), .B0(n113), .C0(n112), .Y(dout[3]) );
  AOI221XL U68 ( .A0(n111), .A1(n75), .B0(n11), .B1(n5), .C0(n110), .Y(n112)
         );
  AOI2BB2XL U69 ( .B0(n102), .B1(n74), .A0N(n115), .A1N(n125), .Y(n113) );
  NAND4BX1 U70 ( .AN(n85), .B(n84), .C(n83), .D(n82), .Y(dout[1]) );
  AOI221XL U71 ( .A0(n9), .A1(n81), .B0(n12), .B1(n7), .C0(n80), .Y(n82) );
  AOI22X1 U72 ( .A0(n8), .A1(n77), .B0(n4), .B1(n76), .Y(n83) );
  CLKINVX3 U73 ( .A(addr[6]), .Y(n6) );
  CLKINVX3 U74 ( .A(n105), .Y(n8) );
  CLKINVX3 U75 ( .A(addr[1]), .Y(n10) );
  CLKINVX3 U76 ( .A(n116), .Y(n14) );
  CLKINVX3 U77 ( .A(n1), .Y(n15) );
  CLKINVX3 U78 ( .A(addr[4]), .Y(n74) );
  CLKINVX3 U79 ( .A(addr[2]), .Y(n75) );
endmodule


module crp_3 ( P, R, K_sub );
  output [1:32] P;
  input [1:32] R;
  input [1:48] K_sub;
  wire   n1;
  wire   [1:48] X;

  sbox1_3 u0 ( .addr(X[1:6]), .dout({P[9], P[17], P[23], P[31]}) );
  sbox2_3 u1 ( .addr({X[7], n1, X[9:12]}), .dout({P[13], P[28], P[2], P[18]})
         );
  sbox3_3 u2 ( .addr(X[13:18]), .dout({P[24], P[16], P[30], P[6]}) );
  sbox4_3 u3 ( .addr(X[19:24]), .dout({P[26], P[20], P[10], P[1]}) );
  sbox5_3 u4 ( .addr(X[25:30]), .dout({P[8], P[14], P[25], P[3]}) );
  sbox6_3 u5 ( .addr(X[31:36]), .dout({P[4], P[29], P[11], P[19]}) );
  sbox7_3 u6 ( .addr(X[37:42]), .dout({P[32], P[12], P[22], P[7]}) );
  sbox8_3 u7 ( .addr(X[43:48]), .dout({P[5], P[27], P[15], P[21]}) );
  XNOR2X1 U1 ( .A(R[5]), .B(K_sub[8]), .Y(X[8]) );
  INVX3 U2 ( .A(X[8]), .Y(n1) );
  CLKXOR2X4 U3 ( .A(R[10]), .B(K_sub[15]), .Y(X[15]) );
  XOR2X1 U4 ( .A(R[1]), .B(K_sub[2]), .Y(X[2]) );
  CLKXOR2X4 U5 ( .A(R[29]), .B(K_sub[42]), .Y(X[42]) );
  CLKXOR2X4 U6 ( .A(R[16]), .B(K_sub[25]), .Y(X[25]) );
  CLKXOR2X4 U7 ( .A(R[8]), .B(K_sub[11]), .Y(X[11]) );
  CLKXOR2X4 U8 ( .A(R[20]), .B(K_sub[31]), .Y(X[31]) );
  CLKXOR2X4 U9 ( .A(R[29]), .B(K_sub[44]), .Y(X[44]) );
  CLKXOR2X4 U10 ( .A(R[16]), .B(K_sub[23]), .Y(X[23]) );
  CLKXOR2X4 U11 ( .A(R[31]), .B(K_sub[46]), .Y(X[46]) );
  CLKXOR2X4 U12 ( .A(R[22]), .B(K_sub[33]), .Y(X[33]) );
  CLKXOR2X4 U13 ( .A(R[12]), .B(K_sub[19]), .Y(X[19]) );
  CLKXOR2X4 U14 ( .A(R[26]), .B(K_sub[39]), .Y(X[39]) );
  CLKXOR2X4 U15 ( .A(R[20]), .B(K_sub[29]), .Y(X[29]) );
  CLKXOR2X2 U16 ( .A(R[4]), .B(K_sub[5]), .Y(X[5]) );
  CLKXOR2X2 U17 ( .A(R[15]), .B(K_sub[22]), .Y(X[22]) );
  CLKXOR2X2 U18 ( .A(R[24]), .B(K_sub[35]), .Y(X[35]) );
  CLKXOR2X2 U19 ( .A(R[21]), .B(K_sub[30]), .Y(X[30]) );
  CLKXOR2X2 U20 ( .A(R[12]), .B(K_sub[17]), .Y(X[17]) );
  CLKXOR2X2 U21 ( .A(R[32]), .B(K_sub[1]), .Y(X[1]) );
  CLKXOR2X2 U22 ( .A(R[13]), .B(K_sub[20]), .Y(X[20]) );
  CLKXOR2X2 U23 ( .A(R[18]), .B(K_sub[27]), .Y(X[27]) );
  CLKXOR2X2 U24 ( .A(R[8]), .B(K_sub[13]), .Y(X[13]) );
  CLKXOR2X2 U25 ( .A(R[5]), .B(K_sub[6]), .Y(X[6]) );
  CLKXOR2X2 U26 ( .A(R[4]), .B(K_sub[7]), .Y(X[7]) );
  CLKXOR2X2 U27 ( .A(R[24]), .B(K_sub[37]), .Y(X[37]) );
  CLKXOR2X2 U28 ( .A(R[28]), .B(K_sub[43]), .Y(X[43]) );
  CLKXOR2X2 U29 ( .A(R[1]), .B(K_sub[48]), .Y(X[48]) );
  CLKXOR2X2 U30 ( .A(R[17]), .B(K_sub[24]), .Y(X[24]) );
  CLKXOR2X2 U31 ( .A(R[9]), .B(K_sub[12]), .Y(X[12]) );
  CLKXOR2X2 U32 ( .A(R[13]), .B(K_sub[18]), .Y(X[18]) );
  CLKXOR2X2 U33 ( .A(R[25]), .B(K_sub[36]), .Y(X[36]) );
  XOR2X1 U34 ( .A(R[23]), .B(K_sub[34]), .Y(X[34]) );
  XOR2X1 U35 ( .A(R[9]), .B(K_sub[14]), .Y(X[14]) );
  XOR2X1 U36 ( .A(R[30]), .B(K_sub[45]), .Y(X[45]) );
  XOR2X1 U37 ( .A(R[21]), .B(K_sub[32]), .Y(X[32]) );
  XOR2X1 U38 ( .A(R[25]), .B(K_sub[38]), .Y(X[38]) );
  XOR2X1 U39 ( .A(R[27]), .B(K_sub[40]), .Y(X[40]) );
  XOR2X1 U40 ( .A(R[3]), .B(K_sub[4]), .Y(X[4]) );
  XOR2X1 U41 ( .A(R[11]), .B(K_sub[16]), .Y(X[16]) );
  XOR2X1 U42 ( .A(R[7]), .B(K_sub[10]), .Y(X[10]) );
  XOR2X1 U43 ( .A(R[14]), .B(K_sub[21]), .Y(X[21]) );
  XOR2X1 U44 ( .A(R[6]), .B(K_sub[9]), .Y(X[9]) );
  XOR2X1 U45 ( .A(R[2]), .B(K_sub[3]), .Y(X[3]) );
  XOR2X1 U46 ( .A(R[28]), .B(K_sub[41]), .Y(X[41]) );
  XOR2X1 U47 ( .A(R[17]), .B(K_sub[26]), .Y(X[26]) );
  XOR2X1 U48 ( .A(R[32]), .B(K_sub[47]), .Y(X[47]) );
  XOR2X1 U49 ( .A(R[19]), .B(K_sub[28]), .Y(X[28]) );
endmodule


module sbox1_2 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127;

  OAI222X4 U13 ( .A0(addr[5]), .A1(n101), .B0(n1), .B1(n100), .C0(n99), .C1(
        n12), .Y(dout[3]) );
  OAI21X2 U42 ( .A0(n4), .A1(n112), .B0(n106), .Y(n123) );
  NAND2X2 U44 ( .A(addr[6]), .B(n8), .Y(n115) );
  NAND2X2 U48 ( .A(addr[1]), .B(n13), .Y(n114) );
  OAI22X2 U49 ( .A0(n69), .A1(n72), .B0(addr[5]), .B1(n120), .Y(n85) );
  NAND2X2 U50 ( .A(n3), .B(n69), .Y(n120) );
  NOR2X2 U51 ( .A(n69), .B(n3), .Y(n124) );
  NOR2X2 U56 ( .A(n109), .B(n3), .Y(n93) );
  NAND2X2 U57 ( .A(addr[1]), .B(addr[6]), .Y(n109) );
  NAND2X2 U59 ( .A(n8), .B(n13), .Y(n112) );
  NOR2X1 U1 ( .A(n114), .B(n120), .Y(n104) );
  AOI221X4 U2 ( .A0(n7), .A1(n90), .B0(n4), .B1(n93), .C0(n102), .Y(n79) );
  NOR3X1 U3 ( .A(n2), .B(addr[6]), .C(n12), .Y(n102) );
  BUFX4 U4 ( .A(addr[4]), .Y(n2) );
  CLKBUFX3 U5 ( .A(addr[2]), .Y(n1) );
  OAI32X1 U6 ( .A0(n112), .A1(n2), .A2(n4), .B0(n115), .B1(n113), .Y(n80) );
  NOR2BXL U7 ( .AN(n118), .B(n1), .Y(n122) );
  CLKBUFX3 U8 ( .A(addr[2]), .Y(n4) );
  OAI221X4 U9 ( .A0(n88), .A1(n72), .B0(addr[5]), .B1(n87), .C0(n86), .Y(
        dout[2]) );
  OAI221X4 U10 ( .A0(addr[5]), .A1(n127), .B0(n126), .B1(n72), .C0(n125), .Y(
        dout[4]) );
  OA21XL U11 ( .A0(n95), .A1(n115), .B0(n107), .Y(n119) );
  AOI222XL U12 ( .A0(n7), .A1(n1), .B0(n2), .B1(n110), .C0(n9), .C1(n12), .Y(
        n111) );
  AOI2BB2X1 U14 ( .B0(n2), .B1(n9), .A0N(addr[4]), .A1N(n115), .Y(n91) );
  BUFX4 U15 ( .A(addr[3]), .Y(n3) );
  CLKINVX1 U16 ( .A(n112), .Y(n7) );
  CLKINVX1 U17 ( .A(n113), .Y(n11) );
  NAND2BX1 U18 ( .AN(n104), .B(n119), .Y(n84) );
  CLKXOR2X2 U19 ( .A(n70), .B(n12), .Y(n90) );
  NOR2X1 U20 ( .A(n69), .B(n70), .Y(n118) );
  OAI21XL U21 ( .A0(n70), .A1(n114), .B0(n91), .Y(n92) );
  NAND2X1 U22 ( .A(n93), .B(n69), .Y(n107) );
  NAND2X1 U23 ( .A(n12), .B(n70), .Y(n113) );
  OAI211X1 U24 ( .A0(n69), .A1(n114), .B0(n108), .C0(n107), .Y(n89) );
  CLKINVX1 U25 ( .A(n109), .Y(n9) );
  NAND2X1 U26 ( .A(n124), .B(n6), .Y(n108) );
  CLKINVX1 U27 ( .A(n114), .Y(n10) );
  CLKINVX1 U28 ( .A(n115), .Y(n6) );
  CLKINVX1 U29 ( .A(n95), .Y(n71) );
  AO22X1 U30 ( .A0(n90), .A1(n6), .B0(n70), .B1(n123), .Y(n76) );
  OAI31X1 U31 ( .A0(n12), .A1(n3), .A2(n8), .B0(n103), .Y(n105) );
  AOI31XL U32 ( .A0(n8), .A1(n12), .A2(n2), .B0(n102), .Y(n103) );
  CLKINVX1 U33 ( .A(addr[6]), .Y(n13) );
  AOI211X1 U34 ( .A0(n5), .A1(n4), .B0(n117), .C0(n116), .Y(n126) );
  CLKINVX1 U35 ( .A(n108), .Y(n5) );
  AOI211X1 U36 ( .A0(n115), .A1(n114), .B0(n113), .C0(n2), .Y(n116) );
  OAI22X1 U37 ( .A0(n120), .A1(n112), .B0(n111), .B1(n70), .Y(n117) );
  AOI211X1 U38 ( .A0(n9), .A1(n118), .B0(n81), .C0(n80), .Y(n88) );
  OAI22X1 U39 ( .A0(n91), .A1(n12), .B0(n3), .B1(n106), .Y(n81) );
  CLKINVX3 U40 ( .A(addr[5]), .Y(n72) );
  NAND2X1 U41 ( .A(n3), .B(n72), .Y(n95) );
  NAND2X1 U43 ( .A(n10), .B(n1), .Y(n106) );
  XOR2X1 U45 ( .A(n82), .B(n2), .Y(n83) );
  NAND2X1 U46 ( .A(n1), .B(n3), .Y(n82) );
  OAI22XL U47 ( .A0(n3), .A1(n8), .B0(n70), .B1(n112), .Y(n94) );
  AOI211XL U52 ( .A0(n98), .A1(n70), .B0(n97), .C0(n104), .Y(n99) );
  OAI22XL U53 ( .A0(n96), .A1(n69), .B0(n95), .B1(n109), .Y(n97) );
  OAI22XL U54 ( .A0(n13), .A1(n72), .B0(n2), .B1(addr[1]), .Y(n98) );
  AOI221XL U55 ( .A0(n71), .A1(addr[6]), .B0(addr[5]), .B1(n94), .C0(n93), .Y(
        n96) );
  OAI21XL U58 ( .A0(addr[1]), .A1(n120), .B0(n119), .Y(n121) );
  AOI221XL U60 ( .A0(n7), .A1(n118), .B0(n93), .B1(n72), .C0(n75), .Y(n78) );
  OAI31X1 U61 ( .A0(n72), .A1(n2), .A2(n74), .B0(n73), .Y(n75) );
  OA21XL U62 ( .A0(n3), .A1(n13), .B0(n109), .Y(n74) );
  OAI21XL U63 ( .A0(n124), .A1(n85), .B0(n10), .Y(n73) );
  OAI21XL U64 ( .A0(n1), .A1(n8), .B0(n109), .Y(n110) );
  INVX4 U65 ( .A(n4), .Y(n12) );
  AOI222XL U66 ( .A0(n124), .A1(n123), .B0(n122), .B1(addr[6]), .C0(n1), .C1(
        n121), .Y(n125) );
  NOR4BBX1 U67 ( .AN(n107), .BN(n106), .C(n105), .D(n104), .Y(n127) );
  AOI222XL U68 ( .A0(n7), .A1(n90), .B0(n89), .B1(n12), .C0(n123), .C1(n69), 
        .Y(n101) );
  AOI2BB2XL U69 ( .B0(addr[5]), .B1(n92), .A0N(n120), .A1N(addr[1]), .Y(n100)
         );
  AOI32X1 U70 ( .A0(n4), .A1(n85), .A2(n7), .B0(n84), .B1(n12), .Y(n86) );
  AOI222XL U71 ( .A0(n124), .A1(n8), .B0(n83), .B1(addr[1]), .C0(n11), .C1(n13), .Y(n87) );
  OAI221X1 U72 ( .A0(n79), .A1(n72), .B0(n4), .B1(n78), .C0(n77), .Y(dout[1])
         );
  AOI32XL U73 ( .A0(addr[6]), .A1(n85), .A2(n1), .B0(n76), .B1(n72), .Y(n77)
         );
  CLKINVX3 U74 ( .A(addr[1]), .Y(n8) );
  CLKINVX3 U75 ( .A(n2), .Y(n69) );
  CLKINVX3 U76 ( .A(n3), .Y(n70) );
endmodule


module sbox2_2 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147;

  NAND2X2 U55 ( .A(n2), .B(n11), .Y(n136) );
  NAND2X2 U57 ( .A(addr[2]), .B(n9), .Y(n104) );
  NAND2X2 U60 ( .A(addr[5]), .B(addr[2]), .Y(n132) );
  NOR2X2 U61 ( .A(n16), .B(n13), .Y(n101) );
  NAND2X2 U62 ( .A(n15), .B(n82), .Y(n146) );
  NAND2X2 U63 ( .A(n3), .B(n83), .Y(n124) );
  NAND2X2 U64 ( .A(addr[6]), .B(n15), .Y(n122) );
  NAND2X2 U67 ( .A(n3), .B(n2), .Y(n133) );
  AOI222XL U1 ( .A0(n4), .A1(n81), .B0(n88), .B1(n83), .C0(n140), .C1(n13), 
        .Y(n89) );
  CLKINVX1 U2 ( .A(n121), .Y(n16) );
  OAI211X4 U3 ( .A0(n147), .A1(n146), .B0(n145), .C0(n144), .Y(dout[4]) );
  NOR2X1 U4 ( .A(n104), .B(n2), .Y(n141) );
  NOR2X1 U5 ( .A(n124), .B(n2), .Y(n140) );
  CLKBUFX4 U6 ( .A(addr[4]), .Y(n2) );
  CLKINVX1 U7 ( .A(addr[5]), .Y(n1) );
  INVX3 U8 ( .A(addr[5]), .Y(n9) );
  NAND3XL U9 ( .A(n98), .B(n97), .C(n96), .Y(dout[1]) );
  NAND2X1 U10 ( .A(addr[1]), .B(addr[6]), .Y(n121) );
  CLKINVX2 U11 ( .A(addr[1]), .Y(n15) );
  OAI221X1 U12 ( .A0(addr[1]), .A1(n136), .B0(n133), .B1(n15), .C0(n87), .Y(
        n95) );
  NAND2X4 U13 ( .A(addr[1]), .B(n82), .Y(n114) );
  INVX3 U14 ( .A(addr[6]), .Y(n82) );
  NAND2XL U15 ( .A(n102), .B(n11), .Y(n109) );
  AOI211XL U16 ( .A0(n10), .A1(n95), .B0(n94), .C0(n93), .Y(n96) );
  AOI2BB2X1 U17 ( .B0(n9), .B1(n12), .A0N(n104), .A1N(n136), .Y(n117) );
  NOR3BXL U18 ( .AN(n135), .B(n134), .C(n4), .Y(n147) );
  BUFX4 U19 ( .A(addr[3]), .Y(n3) );
  NAND2X1 U20 ( .A(n4), .B(n16), .Y(n113) );
  CLKINVX1 U21 ( .A(n146), .Y(n13) );
  CLKINVX1 U22 ( .A(n115), .Y(n4) );
  CLKINVX1 U23 ( .A(n122), .Y(n14) );
  OAI31X1 U24 ( .A0(n124), .A1(n82), .A2(n9), .B0(n123), .Y(n128) );
  OAI21XL U25 ( .A0(n9), .A1(n15), .B0(n140), .Y(n123) );
  OAI22X1 U26 ( .A0(n122), .A1(n124), .B0(n101), .B1(n132), .Y(n84) );
  INVX1 U27 ( .A(n114), .Y(n81) );
  OAI22X1 U28 ( .A0(n122), .A1(n11), .B0(n5), .B1(n121), .Y(n129) );
  NAND3X1 U29 ( .A(n5), .B(n9), .C(n15), .Y(n111) );
  NAND2X1 U30 ( .A(n11), .B(n5), .Y(n115) );
  OAI21XL U31 ( .A0(n83), .A1(n133), .B0(n135), .Y(n85) );
  OAI22XL U32 ( .A0(n117), .A1(n146), .B0(n116), .B1(n132), .Y(n118) );
  AOI222XL U33 ( .A0(n81), .A1(n115), .B0(n6), .B1(n82), .C0(n4), .C1(n13), 
        .Y(n116) );
  CLKINVX1 U34 ( .A(n104), .Y(n8) );
  OAI2BB2XL U35 ( .B0(n114), .B1(n135), .A0N(n126), .A1N(n6), .Y(n106) );
  OAI21XL U36 ( .A0(n112), .A1(n114), .B0(n111), .Y(n120) );
  OAI21XL U37 ( .A0(n133), .A1(n114), .B0(n113), .Y(n119) );
  CLKINVX1 U38 ( .A(n124), .Y(n12) );
  CLKINVX1 U39 ( .A(n136), .Y(n7) );
  CLKINVX1 U40 ( .A(n133), .Y(n6) );
  CLKINVX1 U41 ( .A(n132), .Y(n10) );
  AOI2BB1X1 U42 ( .A0N(n126), .A1N(n125), .B0(n136), .Y(n127) );
  OAI22XL U43 ( .A0(n104), .A1(n114), .B0(n101), .B1(n132), .Y(n102) );
  AO21XL U44 ( .A0(n83), .A1(n7), .B0(n141), .Y(n86) );
  AO21X1 U45 ( .A0(n11), .A1(n8), .B0(n140), .Y(n142) );
  NAND3X1 U46 ( .A(n83), .B(n5), .C(addr[5]), .Y(n135) );
  OAI22X1 U47 ( .A0(addr[5]), .A1(n121), .B0(n122), .B1(n9), .Y(n126) );
  AOI2BB1X1 U48 ( .A0N(n3), .A1N(n1), .B0(n7), .Y(n112) );
  NOR3X1 U49 ( .A(addr[1]), .B(addr[2]), .C(n9), .Y(n125) );
  AOI2BB1XL U50 ( .A0N(n92), .A1N(n91), .B0(addr[5]), .Y(n93) );
  OAI22XL U51 ( .A0(n117), .A1(n114), .B0(n89), .B1(n1), .Y(n94) );
  OAI31XL U52 ( .A0(n114), .A1(n2), .A2(n11), .B0(n90), .Y(n91) );
  OAI21XL U53 ( .A0(n6), .A1(n12), .B0(n14), .Y(n90) );
  NAND2X1 U54 ( .A(n81), .B(n2), .Y(n137) );
  OAI31XL U56 ( .A0(n101), .A1(n3), .A2(addr[2]), .B0(n113), .Y(n92) );
  OAI211X1 U58 ( .A0(n139), .A1(n9), .B0(n138), .C0(n137), .Y(n143) );
  NAND3X1 U59 ( .A(n5), .B(n9), .C(addr[6]), .Y(n138) );
  AOI2BB2X1 U65 ( .B0(n14), .B1(n11), .A0N(n15), .A1N(n136), .Y(n139) );
  OAI22XL U66 ( .A0(addr[5]), .A1(n133), .B0(n3), .B1(n132), .Y(n134) );
  OAI2BB2XL U68 ( .B0(n112), .B1(n122), .A0N(n1), .A1N(n99), .Y(n100) );
  OAI211X1 U69 ( .A0(n146), .A1(n2), .B0(n137), .C0(n113), .Y(n99) );
  NAND3X1 U70 ( .A(n14), .B(n5), .C(n3), .Y(n87) );
  AOI2BB2XL U71 ( .B0(n3), .B1(n105), .A0N(n137), .A1N(n132), .Y(n108) );
  OAI211XL U72 ( .A0(n104), .A1(n146), .B0(n103), .C0(n111), .Y(n105) );
  NAND3XL U73 ( .A(addr[5]), .B(n5), .C(n16), .Y(n103) );
  OAI22XL U74 ( .A0(n3), .A1(n114), .B0(n82), .B1(n115), .Y(n88) );
  NAND4X1 U75 ( .A(n110), .B(n109), .C(n108), .D(n107), .Y(dout[2]) );
  AOI32XL U76 ( .A0(addr[1]), .A1(addr[2]), .A2(n7), .B0(n100), .B1(n83), .Y(
        n110) );
  AOI221XL U77 ( .A0(n125), .A1(addr[4]), .B0(n141), .B1(n14), .C0(n106), .Y(
        n107) );
  AOI33XL U78 ( .A0(n14), .A1(n8), .A2(n2), .B0(n10), .B1(n146), .B2(n3), .Y(
        n145) );
  AOI222XL U79 ( .A0(n143), .A1(n83), .B0(n16), .B1(n142), .C0(n81), .C1(n141), 
        .Y(n144) );
  AOI32XL U80 ( .A0(n8), .A1(n15), .A2(n4), .B0(n13), .B1(n86), .Y(n97) );
  AOI22X1 U81 ( .A0(n16), .A1(n85), .B0(n2), .B1(n84), .Y(n98) );
  NAND2X1 U82 ( .A(n131), .B(n130), .Y(dout[3]) );
  AOI221XL U83 ( .A0(n120), .A1(n83), .B0(addr[2]), .B1(n119), .C0(n118), .Y(
        n131) );
  AOI211X1 U84 ( .A0(n8), .A1(n129), .B0(n128), .C0(n127), .Y(n130) );
  CLKINVX3 U85 ( .A(n2), .Y(n5) );
  CLKINVX3 U86 ( .A(n3), .Y(n11) );
  CLKINVX3 U87 ( .A(addr[2]), .Y(n83) );
endmodule


module sbox3_2 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133;

  NOR2X2 U35 ( .A(n15), .B(addr[3]), .Y(n108) );
  NOR2X2 U50 ( .A(addr[1]), .B(addr[6]), .Y(n107) );
  NOR2X2 U52 ( .A(n20), .B(n2), .Y(n87) );
  NOR2X2 U56 ( .A(n20), .B(n77), .Y(n94) );
  NOR2X1 U1 ( .A(n15), .B(n20), .Y(n106) );
  OAI221X1 U2 ( .A0(n124), .A1(n15), .B0(n3), .B1(addr[1]), .C0(n13), .Y(n104)
         );
  OAI22XL U3 ( .A0(n2), .A1(n77), .B0(n3), .B1(n14), .Y(n123) );
  BUFX4 U4 ( .A(addr[4]), .Y(n2) );
  CLKBUFX3 U5 ( .A(n77), .Y(n1) );
  OAI33X1 U6 ( .A0(n17), .A1(n125), .A2(n77), .B0(n15), .B1(n94), .B2(n119), 
        .Y(n79) );
  INVX3 U7 ( .A(n3), .Y(n77) );
  NOR2X1 U8 ( .A(n9), .B(n3), .Y(n91) );
  NOR2X1 U9 ( .A(n17), .B(n3), .Y(n121) );
  NOR2X1 U10 ( .A(n13), .B(n3), .Y(n95) );
  NOR2X1 U11 ( .A(n3), .B(n2), .Y(n110) );
  CLKBUFX4 U12 ( .A(addr[2]), .Y(n3) );
  OAI221X1 U13 ( .A0(addr[5]), .A1(n90), .B0(n89), .B1(n78), .C0(n88), .Y(
        dout[1]) );
  NOR2X4 U14 ( .A(n10), .B(n76), .Y(n124) );
  NOR2X4 U15 ( .A(addr[3]), .B(n2), .Y(n130) );
  NOR2X4 U16 ( .A(n76), .B(addr[6]), .Y(n125) );
  INVX3 U17 ( .A(addr[1]), .Y(n76) );
  NAND2XL U18 ( .A(n94), .B(n124), .Y(n132) );
  OAI211XL U19 ( .A0(n2), .A1(n8), .B0(n128), .C0(n127), .Y(n129) );
  NAND4XL U20 ( .A(n114), .B(n113), .C(n112), .D(n111), .Y(n115) );
  CLKINVX1 U21 ( .A(n132), .Y(n6) );
  INVX1 U22 ( .A(n124), .Y(n4) );
  CLKINVX1 U23 ( .A(n106), .Y(n14) );
  NAND2X1 U24 ( .A(n9), .B(n11), .Y(n122) );
  CLKINVX1 U25 ( .A(n86), .Y(n11) );
  CLKINVX1 U26 ( .A(n120), .Y(n19) );
  CLKINVX1 U27 ( .A(n119), .Y(n5) );
  CLKINVX1 U28 ( .A(n114), .Y(n7) );
  CLKINVX1 U29 ( .A(n107), .Y(n13) );
  NOR2X1 U30 ( .A(n9), .B(n77), .Y(n103) );
  NOR2X1 U31 ( .A(n4), .B(n77), .Y(n109) );
  INVX1 U32 ( .A(n125), .Y(n12) );
  AOI21X1 U33 ( .A0(n20), .A1(n77), .B0(n94), .Y(n120) );
  OAI21XL U34 ( .A0(n110), .A1(n130), .B0(n124), .Y(n82) );
  CLKINVX1 U36 ( .A(n81), .Y(n9) );
  NOR2X1 U37 ( .A(n12), .B(n15), .Y(n86) );
  NOR2X1 U38 ( .A(n124), .B(n107), .Y(n119) );
  OAI21XL U39 ( .A0(n109), .A1(n91), .B0(n130), .Y(n100) );
  NAND2X1 U40 ( .A(n103), .B(n87), .Y(n114) );
  CLKINVX1 U41 ( .A(n87), .Y(n17) );
  CLKINVX1 U42 ( .A(n91), .Y(n8) );
  CLKINVX1 U43 ( .A(n110), .Y(n18) );
  CLKINVX1 U44 ( .A(n121), .Y(n16) );
  OR2X1 U45 ( .A(n103), .B(n95), .Y(n126) );
  OAI221X1 U46 ( .A0(n12), .A1(n18), .B0(n77), .B1(n11), .C0(n93), .Y(n98) );
  AOI221XL U47 ( .A0(n95), .A1(n2), .B0(n92), .B1(n15), .C0(n6), .Y(n93) );
  OAI21XL U48 ( .A0(n1), .A1(n13), .B0(n8), .Y(n92) );
  XNOR2X1 U49 ( .A(addr[5]), .B(addr[3]), .Y(n102) );
  CLKINVX1 U51 ( .A(addr[5]), .Y(n78) );
  OAI221X1 U53 ( .A0(n13), .A1(n18), .B0(n4), .B1(n17), .C0(n105), .Y(n116) );
  AOI221XL U54 ( .A0(addr[3]), .A1(n104), .B0(n103), .B1(n130), .C0(n6), .Y(
        n105) );
  CLKINVX1 U55 ( .A(addr[6]), .Y(n10) );
  NAND3X1 U57 ( .A(n3), .B(n76), .C(n108), .Y(n113) );
  NOR2X1 U58 ( .A(n10), .B(addr[1]), .Y(n81) );
  AOI32XL U59 ( .A0(n1), .A1(n20), .A2(n124), .B0(n123), .B1(n10), .Y(n128) );
  AOI22XL U60 ( .A0(n2), .A1(n126), .B0(n125), .B1(n130), .Y(n127) );
  AOI222XL U61 ( .A0(n110), .A1(n125), .B0(n109), .B1(n20), .C0(n108), .C1(
        n107), .Y(n111) );
  OAI211XL U62 ( .A0(n106), .A1(n130), .B0(n1), .C0(addr[6]), .Y(n112) );
  OAI21XL U63 ( .A0(n3), .A1(addr[1]), .B0(n12), .Y(n80) );
  AOI221XL U64 ( .A0(n86), .A1(n20), .B0(n87), .B1(n125), .C0(n85), .Y(n89) );
  OAI211X1 U65 ( .A0(n84), .A1(n77), .B0(n83), .C0(n82), .Y(n85) );
  AOI222XL U66 ( .A0(n81), .A1(n20), .B0(n107), .B1(n106), .C0(n130), .C1(n76), 
        .Y(n84) );
  OAI21XL U67 ( .A0(n91), .A1(n6), .B0(addr[4]), .Y(n83) );
  AOI221XL U68 ( .A0(n125), .A1(n19), .B0(addr[3]), .B1(n126), .C0(n96), .Y(
        n97) );
  OAI22X1 U69 ( .A0(n4), .A1(n16), .B0(n14), .B1(n9), .Y(n96) );
  OAI211X1 U70 ( .A0(n13), .A1(n16), .B0(n118), .C0(n117), .Y(dout[3]) );
  AOI32XL U71 ( .A0(n125), .A1(n3), .A2(n102), .B0(n108), .B1(n109), .Y(n118)
         );
  AOI22XL U72 ( .A0(n116), .A1(n78), .B0(addr[5]), .B1(n115), .Y(n117) );
  AOI221XL U73 ( .A0(n121), .A1(n125), .B0(n95), .B1(n108), .C0(n7), .Y(n88)
         );
  AOI221XL U74 ( .A0(n130), .A1(n80), .B0(n94), .B1(n122), .C0(n79), .Y(n90)
         );
  NAND4X1 U75 ( .A(n101), .B(n113), .C(n100), .D(n99), .Y(dout[2]) );
  NAND3XL U76 ( .A(n2), .B(n124), .C(n102), .Y(n101) );
  AOI2BB2XL U77 ( .B0(addr[5]), .B1(n98), .A0N(addr[5]), .A1N(n97), .Y(n99) );
  OAI221X1 U78 ( .A0(n133), .A1(n78), .B0(n2), .B1(n132), .C0(n131), .Y(
        dout[4]) );
  AOI32XL U79 ( .A0(n130), .A1(n10), .A2(addr[2]), .B0(n129), .B1(n78), .Y(
        n131) );
  AOI222XL U80 ( .A0(n19), .A1(n122), .B0(n121), .B1(addr[1]), .C0(n120), .C1(
        n5), .Y(n133) );
  CLKINVX3 U81 ( .A(n2), .Y(n15) );
  CLKINVX3 U82 ( .A(addr[3]), .Y(n20) );
endmodule


module sbox4_2 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126;

  OAI32X4 U12 ( .A0(n12), .A1(n2), .A2(addr[2]), .B0(n11), .B1(n108), .Y(n123)
         );
  OAI222X4 U20 ( .A0(addr[2]), .A1(n92), .B0(n106), .B1(n91), .C0(n90), .C1(
        n14), .Y(dout[2]) );
  OAI222X4 U33 ( .A0(addr[4]), .A1(n106), .B0(n6), .B1(n108), .C0(n2), .C1(
        n118), .Y(n83) );
  NAND2X2 U34 ( .A(addr[4]), .B(n2), .Y(n108) );
  NOR2X2 U43 ( .A(n72), .B(addr[4]), .Y(n113) );
  NOR2X2 U45 ( .A(n11), .B(n2), .Y(n111) );
  NAND2X2 U51 ( .A(n6), .B(n71), .Y(n118) );
  NOR2X2 U52 ( .A(n16), .B(addr[5]), .Y(n97) );
  NAND2X2 U53 ( .A(addr[6]), .B(addr[1]), .Y(n85) );
  NAND2X2 U54 ( .A(addr[1]), .B(n71), .Y(n116) );
  NOR2X2 U55 ( .A(n115), .B(n11), .Y(n121) );
  NAND2X2 U56 ( .A(n72), .B(n16), .Y(n115) );
  NAND2X2 U57 ( .A(addr[5]), .B(n16), .Y(n96) );
  NAND2X2 U58 ( .A(addr[6]), .B(n6), .Y(n106) );
  OAI222X1 U1 ( .A0(n12), .A1(n85), .B0(n97), .B1(n116), .C0(n16), .C1(n118), 
        .Y(n73) );
  CLKINVX1 U2 ( .A(n116), .Y(n9) );
  OAI31X4 U3 ( .A0(n118), .A1(n11), .A2(n16), .B0(n117), .Y(n119) );
  CLKINVX1 U4 ( .A(n72), .Y(n1) );
  CLKBUFX3 U5 ( .A(addr[3]), .Y(n2) );
  OAI221X1 U6 ( .A0(addr[2]), .A1(n80), .B0(n118), .B1(n105), .C0(n79), .Y(
        dout[1]) );
  INVX4 U7 ( .A(addr[5]), .Y(n11) );
  OAI31X1 U8 ( .A0(n108), .A1(addr[5]), .A2(n5), .B0(n107), .Y(n109) );
  AOI222XL U9 ( .A0(n16), .A1(n71), .B0(n113), .B1(n6), .C0(addr[1]), .C1(n72), 
        .Y(n114) );
  OAI222X1 U10 ( .A0(addr[1]), .A1(n84), .B0(n85), .B1(n74), .C0(n72), .C1(
        n107), .Y(n75) );
  NAND2XL U11 ( .A(n1), .B(addr[5]), .Y(n84) );
  AOI211XL U13 ( .A0(n83), .A1(n11), .B0(n82), .C0(n7), .Y(n92) );
  NAND2XL U14 ( .A(n16), .B(n11), .Y(n74) );
  CLKINVX1 U15 ( .A(n118), .Y(n3) );
  CLKINVX1 U16 ( .A(n115), .Y(n15) );
  CLKINVX1 U17 ( .A(n112), .Y(n4) );
  OAI21X1 U18 ( .A0(n9), .A1(n5), .B0(n14), .Y(n112) );
  AOI22X1 U19 ( .A0(n10), .A1(n111), .B0(n5), .B1(n113), .Y(n93) );
  OAI211X1 U21 ( .A0(n6), .A1(n115), .B0(n93), .C0(n8), .Y(n94) );
  CLKINVX1 U22 ( .A(n85), .Y(n10) );
  NAND2X1 U23 ( .A(n97), .B(n72), .Y(n105) );
  NAND2X1 U24 ( .A(n113), .B(n3), .Y(n98) );
  NAND2X1 U25 ( .A(n9), .B(n97), .Y(n107) );
  NAND2X1 U26 ( .A(n118), .B(n85), .Y(n110) );
  OAI21XL U27 ( .A0(n15), .A1(n11), .B0(n108), .Y(n95) );
  CLKINVX1 U28 ( .A(n84), .Y(n13) );
  CLKINVX1 U29 ( .A(addr[2]), .Y(n14) );
  OAI31X1 U30 ( .A0(n16), .A1(addr[6]), .A2(n11), .B0(n87), .Y(n88) );
  OAI21XL U31 ( .A0(n113), .A1(n12), .B0(n10), .Y(n87) );
  OAI211X1 U32 ( .A0(n76), .A1(n16), .B0(n98), .C0(n8), .Y(n77) );
  AOI222XL U35 ( .A0(addr[5]), .A1(addr[6]), .B0(n111), .B1(addr[1]), .C0(n5), 
        .C1(n2), .Y(n76) );
  NAND3XL U36 ( .A(n10), .B(n72), .C(addr[4]), .Y(n117) );
  OAI22XL U37 ( .A0(n116), .A1(n115), .B0(n1), .B1(n112), .Y(n78) );
  CLKINVX3 U38 ( .A(addr[4]), .Y(n16) );
  OAI2BB2XL U39 ( .B0(n115), .B1(n106), .A0N(n11), .A1N(n86), .Y(n89) );
  OAI221XL U40 ( .A0(n116), .A1(addr[4]), .B0(n108), .B1(addr[1]), .C0(n117), 
        .Y(n86) );
  CLKINVX1 U41 ( .A(addr[6]), .Y(n71) );
  CLKINVX1 U42 ( .A(n81), .Y(n7) );
  OAI21XL U44 ( .A0(n96), .A1(n118), .B0(n93), .Y(n82) );
  NAND3X1 U46 ( .A(n101), .B(n100), .C(n99), .Y(n102) );
  AOI32X1 U47 ( .A0(n96), .A1(n72), .A2(n9), .B0(n10), .B1(n95), .Y(n101) );
  AOI2BB2XL U48 ( .B0(n6), .B1(n121), .A0N(n98), .A1N(addr[5]), .Y(n99) );
  OAI21XL U49 ( .A0(n97), .A1(n12), .B0(n5), .Y(n100) );
  AOI2BB2XL U50 ( .B0(n5), .B1(n123), .A0N(n122), .A1N(n14), .Y(n124) );
  AOI211XL U59 ( .A0(n5), .A1(n121), .B0(n120), .C0(n119), .Y(n122) );
  OAI22XL U60 ( .A0(n116), .A1(n115), .B0(addr[5]), .B1(n114), .Y(n120) );
  CLKINVX1 U61 ( .A(n75), .Y(n8) );
  AOI32XL U62 ( .A0(n9), .A1(n96), .A2(n1), .B0(addr[1]), .B1(n121), .Y(n81)
         );
  AOI222XL U63 ( .A0(n5), .A1(n12), .B0(n121), .B1(n116), .C0(n2), .C1(n73), 
        .Y(n80) );
  AOI22XL U64 ( .A0(n78), .A1(n11), .B0(addr[2]), .B1(n77), .Y(n79) );
  NAND2XL U65 ( .A(n111), .B(addr[4]), .Y(n91) );
  AOI211X1 U66 ( .A0(n13), .A1(n110), .B0(n89), .C0(n88), .Y(n90) );
  OAI211X1 U67 ( .A0(n106), .A1(n105), .B0(n104), .C0(n103), .Y(dout[3]) );
  AOI32X1 U68 ( .A0(n2), .A1(n12), .A2(n9), .B0(n94), .B1(n14), .Y(n104) );
  AOI22XL U69 ( .A0(addr[2]), .A1(n102), .B0(n3), .B1(n123), .Y(n103) );
  OAI211X1 U70 ( .A0(addr[2]), .A1(n126), .B0(n125), .C0(n124), .Y(dout[4]) );
  AOI32X1 U71 ( .A0(n10), .A1(n12), .A2(n2), .B0(n4), .B1(n13), .Y(n125) );
  AOI221XL U72 ( .A0(n3), .A1(n111), .B0(n15), .B1(n110), .C0(n109), .Y(n126)
         );
  CLKINVX3 U73 ( .A(n106), .Y(n5) );
  CLKINVX3 U74 ( .A(addr[1]), .Y(n6) );
  CLKINVX3 U75 ( .A(n96), .Y(n12) );
  CLKINVX3 U76 ( .A(n2), .Y(n72) );
endmodule


module sbox5_2 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121;

  OAI222X4 U18 ( .A0(addr[3]), .A1(n106), .B0(n68), .B1(n90), .C0(n6), .C1(n13), .Y(n93) );
  OAI22X2 U40 ( .A0(addr[5]), .A1(n106), .B0(n69), .B1(n114), .Y(n116) );
  NOR2X2 U41 ( .A(n3), .B(addr[3]), .Y(n102) );
  NAND2X2 U45 ( .A(addr[6]), .B(n13), .Y(n114) );
  NAND2X2 U50 ( .A(n13), .B(n68), .Y(n110) );
  NAND2X2 U52 ( .A(addr[1]), .B(n68), .Y(n113) );
  NAND2X2 U54 ( .A(addr[1]), .B(addr[6]), .Y(n106) );
  NAND2X2 U55 ( .A(addr[3]), .B(n6), .Y(n121) );
  CLKINVX1 U1 ( .A(addr[5]), .Y(n1) );
  AOI221XL U2 ( .A0(n93), .A1(n1), .B0(n14), .B1(n8), .C0(n92), .Y(n105) );
  INVX3 U3 ( .A(addr[5]), .Y(n69) );
  OAI221X4 U4 ( .A0(n111), .A1(n110), .B0(n121), .B1(n114), .C0(n109), .Y(n112) );
  OAI221X4 U5 ( .A0(n6), .A1(n114), .B0(n69), .B1(n113), .C0(n120), .Y(n115)
         );
  OAI221X4 U6 ( .A0(n107), .A1(n121), .B0(n111), .B1(n113), .C0(n85), .Y(n86)
         );
  OAI31X1 U7 ( .A0(n70), .A1(addr[5]), .A2(addr[1]), .B0(n81), .Y(n73) );
  OAI32X1 U8 ( .A0(n114), .A1(addr[5]), .A2(n3), .B0(n5), .B1(n107), .Y(n79)
         );
  AOI32XL U9 ( .A0(n8), .A1(n98), .A2(n16), .B0(n2), .B1(n73), .Y(n77) );
  CLKBUFX3 U10 ( .A(addr[4]), .Y(n2) );
  CLKINVX1 U11 ( .A(n81), .Y(n7) );
  NAND2X1 U12 ( .A(n10), .B(n8), .Y(n81) );
  CLKINVX1 U13 ( .A(n110), .Y(n12) );
  CLKXOR2X2 U14 ( .A(n70), .B(n69), .Y(n94) );
  AOI2BB1X1 U15 ( .A0N(n6), .A1N(n1), .B0(n8), .Y(n111) );
  NOR2X1 U16 ( .A(n121), .B(n69), .Y(n91) );
  NOR2BX1 U17 ( .AN(n116), .B(n90), .Y(n83) );
  NAND2X1 U19 ( .A(n12), .B(n69), .Y(n120) );
  CLKINVX1 U20 ( .A(n113), .Y(n16) );
  NAND2X1 U21 ( .A(n16), .B(n69), .Y(n107) );
  CLKINVX1 U22 ( .A(n121), .Y(n5) );
  OAI31X1 U23 ( .A0(n4), .A1(n8), .A2(n113), .B0(n99), .Y(n72) );
  CLKINVX1 U24 ( .A(n106), .Y(n14) );
  OAI2BB2XL U25 ( .B0(n1), .B1(n113), .A0N(n98), .A1N(n10), .Y(n101) );
  CLKINVX1 U26 ( .A(n114), .Y(n10) );
  CLKINVX1 U27 ( .A(n90), .Y(n9) );
  CLKINVX1 U28 ( .A(addr[1]), .Y(n13) );
  CLKINVX1 U29 ( .A(addr[3]), .Y(n70) );
  CLKINVX1 U30 ( .A(addr[6]), .Y(n68) );
  AOI211X1 U31 ( .A0(n91), .A1(addr[1]), .B0(n80), .C0(n79), .Y(n89) );
  OAI2BB2XL U32 ( .B0(n111), .B1(n106), .A0N(n94), .A1N(n12), .Y(n80) );
  AOI211X1 U33 ( .A0(n102), .A1(n84), .B0(n83), .C0(n82), .Y(n85) );
  OAI21XL U34 ( .A0(n68), .A1(n1), .B0(n106), .Y(n84) );
  NOR3XL U35 ( .A(n94), .B(n3), .C(n110), .Y(n82) );
  AOI222XL U36 ( .A0(n14), .A1(n9), .B0(addr[5]), .B1(n108), .C0(n15), .C1(n6), 
        .Y(n109) );
  CLKINVX1 U37 ( .A(n107), .Y(n15) );
  OAI21XL U38 ( .A0(addr[6]), .A1(addr[3]), .B0(n106), .Y(n108) );
  NAND2X1 U39 ( .A(addr[3]), .B(n3), .Y(n90) );
  NAND2X1 U42 ( .A(n2), .B(addr[5]), .Y(n98) );
  NAND2X1 U43 ( .A(n3), .B(n70), .Y(n97) );
  OAI21XL U44 ( .A0(addr[1]), .A1(n97), .B0(n96), .Y(n103) );
  AOI33XL U46 ( .A0(n3), .A1(n95), .A2(addr[5]), .B0(n94), .B1(n6), .B2(
        addr[1]), .Y(n96) );
  OAI21XL U47 ( .A0(n13), .A1(n70), .B0(n114), .Y(n95) );
  OAI21XL U48 ( .A0(addr[6]), .A1(n121), .B0(n99), .Y(n100) );
  NAND2X1 U49 ( .A(n71), .B(n12), .Y(n99) );
  XOR2X1 U51 ( .A(n4), .B(n3), .Y(n71) );
  AOI2BB2XL U53 ( .B0(n102), .B1(n116), .A0N(n2), .A1N(n75), .Y(n76) );
  AOI211X1 U56 ( .A0(n11), .A1(n3), .B0(n74), .C0(n83), .Y(n75) );
  AO22XL U57 ( .A0(n16), .A1(n5), .B0(addr[6]), .B1(n102), .Y(n74) );
  CLKINVX1 U58 ( .A(n120), .Y(n11) );
  CLKINVX1 U59 ( .A(n2), .Y(n4) );
  AO22XL U60 ( .A0(n16), .A1(n9), .B0(addr[6]), .B1(n91), .Y(n92) );
  AOI222XL U61 ( .A0(n116), .A1(n6), .B0(addr[3]), .B1(n115), .C0(n16), .C1(n8), .Y(n117) );
  OAI221X1 U62 ( .A0(n2), .A1(n105), .B0(n110), .B1(n121), .C0(n104), .Y(
        dout[3]) );
  AOI222XL U63 ( .A0(n2), .A1(n103), .B0(n102), .B1(n101), .C0(n100), .C1(n1), 
        .Y(n104) );
  OAI211X1 U64 ( .A0(n2), .A1(n89), .B0(n88), .C0(n87), .Y(dout[2]) );
  AOI33XL U65 ( .A0(n5), .A1(n98), .A2(n10), .B0(n3), .B1(n94), .B2(n12), .Y(
        n88) );
  AOI222XL U66 ( .A0(n7), .A1(n69), .B0(n2), .B1(n86), .C0(n91), .C1(n14), .Y(
        n87) );
  OAI211X1 U67 ( .A0(n78), .A1(n69), .B0(n77), .C0(n76), .Y(dout[1]) );
  AOI221XL U68 ( .A0(n5), .A1(addr[1]), .B0(n14), .B1(n8), .C0(n72), .Y(n78)
         );
  OAI211X1 U69 ( .A0(n121), .A1(n120), .B0(n119), .C0(n118), .Y(dout[4]) );
  AOI32XL U70 ( .A0(n8), .A1(n114), .A2(addr[5]), .B0(n2), .B1(n112), .Y(n119)
         );
  AOI2BB2X1 U71 ( .B0(n7), .B1(n69), .A0N(n2), .A1N(n117), .Y(n118) );
  BUFX4 U72 ( .A(addr[2]), .Y(n3) );
  CLKINVX3 U73 ( .A(n3), .Y(n6) );
  CLKINVX3 U74 ( .A(n97), .Y(n8) );
endmodule


module sbox6_2 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147;

  NAND2X2 U39 ( .A(n138), .B(addr[3]), .Y(n147) );
  NOR2X2 U47 ( .A(n84), .B(n82), .Y(n138) );
  NOR2X2 U50 ( .A(n14), .B(n4), .Y(n119) );
  NOR2X2 U58 ( .A(n9), .B(n14), .Y(n125) );
  NAND2X2 U61 ( .A(n97), .B(n103), .Y(n112) );
  NOR2X2 U62 ( .A(n18), .B(addr[1]), .Y(n103) );
  NOR2X2 U63 ( .A(n9), .B(addr[3]), .Y(n97) );
  NAND2X2 U64 ( .A(n117), .B(n131), .Y(n140) );
  NOR2X2 U65 ( .A(n5), .B(addr[3]), .Y(n131) );
  NOR2X2 U66 ( .A(n85), .B(addr[6]), .Y(n117) );
  NOR2X1 U1 ( .A(n84), .B(addr[3]), .Y(n102) );
  AOI211X1 U2 ( .A0(n13), .A1(n14), .B0(n131), .C0(n143), .Y(n121) );
  CLKINVX1 U3 ( .A(addr[3]), .Y(n1) );
  INVX3 U4 ( .A(addr[3]), .Y(n14) );
  CLKINVX1 U5 ( .A(n9), .Y(n2) );
  INVX4 U6 ( .A(n4), .Y(n9) );
  CLKBUFX3 U7 ( .A(addr[4]), .Y(n4) );
  CLKINVX1 U8 ( .A(n84), .Y(n3) );
  OAI222X1 U9 ( .A0(n91), .A1(n13), .B0(n5), .B1(n8), .C0(addr[5]), .C1(n10), 
        .Y(n92) );
  BUFX4 U10 ( .A(addr[2]), .Y(n5) );
  OAI221X1 U11 ( .A0(n18), .A1(n7), .B0(n14), .B1(n16), .C0(n86), .Y(n90) );
  INVX3 U12 ( .A(n96), .Y(n16) );
  OAI221X4 U13 ( .A0(n123), .A1(n17), .B0(n82), .B1(n13), .C0(n15), .Y(n124)
         );
  NOR2X4 U14 ( .A(addr[1]), .B(addr[6]), .Y(n130) );
  NOR2X4 U15 ( .A(n5), .B(addr[5]), .Y(n143) );
  INVX1 U16 ( .A(n130), .Y(n83) );
  CLKINVX1 U17 ( .A(n125), .Y(n7) );
  NAND2X1 U18 ( .A(n83), .B(n16), .Y(n105) );
  INVXL U19 ( .A(n121), .Y(n12) );
  CLKINVX1 U20 ( .A(n138), .Y(n81) );
  CLKINVX1 U21 ( .A(n117), .Y(n82) );
  CLKINVX1 U22 ( .A(n119), .Y(n10) );
  NOR2X1 U23 ( .A(n16), .B(n123), .Y(n144) );
  NOR2X1 U24 ( .A(n85), .B(n18), .Y(n96) );
  CLKINVX1 U25 ( .A(n103), .Y(n17) );
  OAI211X1 U26 ( .A0(n83), .A1(n7), .B0(n104), .C0(n112), .Y(n108) );
  OAI21XL U27 ( .A0(n103), .A1(n117), .B0(n102), .Y(n104) );
  OAI21XL U28 ( .A0(n132), .A1(n18), .B0(n1), .Y(n86) );
  AOI21X1 U29 ( .A0(n9), .A1(n102), .B0(n125), .Y(n91) );
  OAI2BB2XL U30 ( .B0(n143), .B1(n83), .A0N(n143), .A1N(n117), .Y(n118) );
  CLKINVX1 U31 ( .A(n122), .Y(n15) );
  CLKINVX1 U32 ( .A(n126), .Y(n11) );
  CLKINVX1 U33 ( .A(n97), .Y(n8) );
  NAND2BX1 U34 ( .AN(n144), .B(n137), .Y(n107) );
  CLKINVX1 U35 ( .A(addr[1]), .Y(n85) );
  NOR2X1 U36 ( .A(n16), .B(n3), .Y(n122) );
  NOR2X1 U37 ( .A(addr[1]), .B(n2), .Y(n132) );
  OAI22X1 U38 ( .A0(n10), .A1(n82), .B0(n5), .B1(n11), .Y(n88) );
  NAND2X1 U40 ( .A(n3), .B(n13), .Y(n123) );
  NAND4X1 U41 ( .A(n147), .B(n140), .C(n100), .D(n99), .Y(n101) );
  AOI222XL U42 ( .A0(n98), .A1(n84), .B0(n102), .B1(n130), .C0(n97), .C1(n105), 
        .Y(n99) );
  NAND3X1 U43 ( .A(n5), .B(n10), .C(n96), .Y(n100) );
  OAI221X1 U44 ( .A0(n14), .A1(n17), .B0(n10), .B1(n18), .C0(n11), .Y(n98) );
  AOI22X1 U45 ( .A0(n4), .A1(n115), .B0(addr[5]), .B1(n114), .Y(n129) );
  OAI21XL U46 ( .A0(n121), .A1(n83), .B0(n147), .Y(n115) );
  OAI21XL U48 ( .A0(n113), .A1(n84), .B0(n112), .Y(n114) );
  AOI221XL U49 ( .A0(n119), .A1(n85), .B0(n130), .B1(addr[3]), .C0(n111), .Y(
        n113) );
  OAI22XL U51 ( .A0(n82), .A1(n9), .B0(addr[3]), .B1(n16), .Y(n111) );
  OAI22XL U52 ( .A0(n14), .A1(n18), .B0(addr[1]), .B1(n10), .Y(n142) );
  AOI211X1 U53 ( .A0(n4), .A1(n135), .B0(n134), .C0(n133), .Y(n136) );
  OA21XL U54 ( .A0(n1), .A1(n3), .B0(n132), .Y(n133) );
  OAI2BB2XL U55 ( .B0(n2), .B1(n15), .A0N(n131), .A1N(n130), .Y(n134) );
  OAI22X1 U56 ( .A0(n5), .A1(n82), .B0(n84), .B1(n16), .Y(n135) );
  CLKINVX3 U57 ( .A(addr[5]), .Y(n13) );
  AOI2BB2X1 U59 ( .B0(n5), .B1(n130), .A0N(n3), .A1N(n17), .Y(n137) );
  NOR2X1 U60 ( .A(n17), .B(n2), .Y(n126) );
  AOI2BB2XL U67 ( .B0(n143), .B1(n90), .A0N(n89), .A1N(n13), .Y(n94) );
  AOI211X1 U68 ( .A0(n122), .A1(n4), .B0(n88), .C0(n87), .Y(n89) );
  OAI32X1 U69 ( .A0(n17), .A1(n14), .A2(n84), .B0(n81), .B1(n8), .Y(n87) );
  NAND3X1 U70 ( .A(n147), .B(n140), .C(n139), .Y(n141) );
  AOI32X1 U71 ( .A0(n5), .A1(n85), .A2(n4), .B0(n138), .B1(n9), .Y(n139) );
  AO22XL U72 ( .A0(n143), .A1(n2), .B0(n116), .B1(n9), .Y(n120) );
  OAI21XL U73 ( .A0(n3), .A1(n13), .B0(n123), .Y(n116) );
  CLKINVX1 U74 ( .A(n106), .Y(n6) );
  AOI32XL U75 ( .A0(n105), .A1(n9), .A2(n1), .B0(addr[1]), .B1(n125), .Y(n106)
         );
  OAI211X1 U76 ( .A0(n9), .A1(n140), .B0(n110), .C0(n109), .Y(dout[2]) );
  AOI222XL U77 ( .A0(n108), .A1(n13), .B0(n143), .B1(n6), .C0(n119), .C1(n107), 
        .Y(n109) );
  AOI2BB2XL U78 ( .B0(addr[5]), .B1(n101), .A0N(n84), .A1N(n112), .Y(n110) );
  OAI211X1 U79 ( .A0(n2), .A1(n147), .B0(n146), .C0(n145), .Y(dout[4]) );
  AOI222XL U80 ( .A0(n144), .A1(n14), .B0(n143), .B1(n142), .C0(n141), .C1(n13), .Y(n145) );
  OA22X1 U81 ( .A0(n7), .A1(n137), .B0(n136), .B1(n13), .Y(n146) );
  NAND3X1 U82 ( .A(n129), .B(n128), .C(n127), .Y(dout[3]) );
  AOI32XL U83 ( .A0(n120), .A1(n14), .A2(addr[1]), .B0(n119), .B1(n118), .Y(
        n128) );
  AOI222XL U84 ( .A0(n144), .A1(n9), .B0(n126), .B1(n12), .C0(n125), .C1(n124), 
        .Y(n127) );
  NAND3BX1 U85 ( .AN(n95), .B(n94), .C(n93), .Y(dout[1]) );
  OAI222X1 U86 ( .A0(n140), .A1(n4), .B0(n112), .B1(n84), .C0(n16), .C1(n91), 
        .Y(n95) );
  AOI32XL U87 ( .A0(addr[1]), .A1(n13), .A2(n125), .B0(n130), .B1(n92), .Y(n93) );
  CLKINVX3 U88 ( .A(addr[6]), .Y(n18) );
  CLKINVX3 U89 ( .A(n5), .Y(n84) );
endmodule


module sbox7_2 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148;

  OAI222X4 U19 ( .A0(n11), .A1(n129), .B0(n4), .B1(n8), .C0(addr[1]), .C1(n21), 
        .Y(n122) );
  OAI33X4 U33 ( .A0(addr[1]), .A1(n4), .A2(n5), .B0(n9), .B1(n85), .B2(n84), 
        .Y(n97) );
  NOR2X2 U44 ( .A(n87), .B(n4), .Y(n116) );
  NOR2X2 U48 ( .A(addr[1]), .B(addr[6]), .Y(n136) );
  NOR2X2 U51 ( .A(n16), .B(n87), .Y(n125) );
  NOR2X2 U52 ( .A(n9), .B(addr[3]), .Y(n131) );
  NOR2X2 U58 ( .A(n93), .B(n124), .Y(n142) );
  NOR2X2 U60 ( .A(n10), .B(addr[1]), .Y(n93) );
  NOR2X2 U62 ( .A(n83), .B(n3), .Y(n137) );
  NOR2X2 U65 ( .A(n10), .B(n86), .Y(n140) );
  NAND2X1 U1 ( .A(n3), .B(n4), .Y(n119) );
  CLKBUFX3 U2 ( .A(addr[4]), .Y(n4) );
  CLKINVX1 U3 ( .A(n83), .Y(n1) );
  CLKINVX1 U4 ( .A(n85), .Y(n2) );
  CLKBUFX3 U5 ( .A(addr[2]), .Y(n5) );
  OAI31X1 U6 ( .A0(n87), .A1(n83), .A2(n86), .B0(n117), .Y(n121) );
  NOR2X4 U7 ( .A(n86), .B(addr[6]), .Y(n124) );
  OAI22X1 U8 ( .A0(addr[1]), .A1(n21), .B0(n5), .B1(n113), .Y(n100) );
  OAI22X1 U9 ( .A0(n4), .A1(n16), .B0(addr[3]), .B1(n19), .Y(n103) );
  AOI211XL U10 ( .A0(n5), .A1(n7), .B0(n131), .C0(n130), .Y(n132) );
  NOR3XL U11 ( .A(n11), .B(addr[3]), .C(n2), .Y(n130) );
  OAI21XL U12 ( .A0(n3), .A1(n1), .B0(n119), .Y(n89) );
  BUFX4 U13 ( .A(addr[5]), .Y(n3) );
  AOI221XL U14 ( .A0(n140), .A1(n89), .B0(n109), .B1(n7), .C0(n88), .Y(n96) );
  CLKINVX1 U15 ( .A(n140), .Y(n9) );
  OAI2BB2XL U16 ( .B0(n142), .B1(n19), .A0N(n141), .A1N(n140), .Y(n143) );
  CLKINVX1 U17 ( .A(n125), .Y(n14) );
  CLKINVX1 U18 ( .A(n142), .Y(n7) );
  NAND2X1 U20 ( .A(n14), .B(n20), .Y(n105) );
  CLKINVX1 U21 ( .A(n123), .Y(n15) );
  CLKINVX1 U22 ( .A(n109), .Y(n18) );
  NAND2X1 U23 ( .A(n124), .B(n87), .Y(n113) );
  CLKINVX1 U24 ( .A(n137), .Y(n19) );
  NOR2X1 U25 ( .A(n19), .B(n87), .Y(n109) );
  CLKINVX1 U26 ( .A(n136), .Y(n11) );
  OAI22XL U27 ( .A0(n137), .A1(n8), .B0(n86), .B1(n18), .Y(n146) );
  OAI21X1 U28 ( .A0(n83), .A1(n14), .B0(n129), .Y(n141) );
  NAND2X1 U29 ( .A(n116), .B(n16), .Y(n129) );
  CLKINVX1 U30 ( .A(n93), .Y(n6) );
  OAI21XL U31 ( .A0(n119), .A1(n6), .B0(n118), .Y(n120) );
  OAI21XL U32 ( .A0(n125), .A1(n137), .B0(n124), .Y(n118) );
  NOR2X1 U34 ( .A(n16), .B(n21), .Y(n123) );
  CLKINVX1 U35 ( .A(n145), .Y(n21) );
  OAI22XL U36 ( .A0(n137), .A1(n113), .B0(n10), .B1(n15), .Y(n88) );
  CLKINVX1 U37 ( .A(n116), .Y(n84) );
  CLKINVX1 U38 ( .A(n131), .Y(n8) );
  CLKINVX1 U39 ( .A(n134), .Y(n20) );
  NOR2XL U40 ( .A(n125), .B(n83), .Y(n110) );
  CLKINVX1 U41 ( .A(n119), .Y(n17) );
  CLKINVX1 U42 ( .A(n103), .Y(n12) );
  OA21XL U43 ( .A0(n13), .A1(n6), .B0(n117), .Y(n102) );
  CLKINVX1 U45 ( .A(n105), .Y(n13) );
  OAI2BB1XL U46 ( .A0N(n103), .A1N(n124), .B0(n102), .Y(n104) );
  OAI22X1 U47 ( .A0(n16), .A1(n84), .B0(n4), .B1(n20), .Y(n112) );
  NOR4X1 U49 ( .A(n4), .B(addr[3]), .C(n86), .D(n85), .Y(n99) );
  XNOR2X1 U50 ( .A(addr[6]), .B(n5), .Y(n101) );
  AOI211X1 U53 ( .A0(n116), .A1(addr[6]), .B0(n115), .C0(n114), .Y(n128) );
  OAI222X1 U54 ( .A0(n111), .A1(n9), .B0(n110), .B1(n6), .C0(n11), .C1(n18), 
        .Y(n115) );
  OAI2BB2XL U55 ( .B0(n17), .B1(n113), .A0N(n86), .A1N(n112), .Y(n114) );
  OA21XL U56 ( .A0(n87), .A1(n3), .B0(n15), .Y(n111) );
  NAND2X1 U57 ( .A(n5), .B(n136), .Y(n133) );
  CLKINVX1 U59 ( .A(addr[6]), .Y(n10) );
  AOI211X1 U61 ( .A0(n131), .A1(n3), .B0(n92), .C0(n91), .Y(n95) );
  OAI221X1 U63 ( .A0(n86), .A1(n21), .B0(n9), .B1(n19), .C0(n102), .Y(n92) );
  OAI31X1 U64 ( .A0(n87), .A1(n83), .A2(n11), .B0(n90), .Y(n91) );
  AO21XL U66 ( .A0(n119), .A1(n129), .B0(addr[6]), .Y(n90) );
  NOR2X1 U67 ( .A(n83), .B(addr[3]), .Y(n145) );
  AOI21XL U68 ( .A0(addr[3]), .A1(n98), .B0(n97), .Y(n108) );
  OAI2BB1XL U69 ( .A0N(n85), .A1N(n124), .B0(n133), .Y(n98) );
  NAND3X1 U70 ( .A(n136), .B(n87), .C(n3), .Y(n117) );
  NOR2X1 U71 ( .A(addr[3]), .B(n3), .Y(n134) );
  OAI21X1 U72 ( .A0(n5), .A1(n142), .B0(n133), .Y(n138) );
  OAI22XL U73 ( .A0(n142), .A1(n84), .B0(n1), .B1(n132), .Y(n135) );
  AO21X1 U74 ( .A0(n139), .A1(n16), .B0(n138), .Y(n144) );
  OAI21XL U75 ( .A0(n2), .A1(n86), .B0(n6), .Y(n139) );
  OAI221X1 U76 ( .A0(n96), .A1(n85), .B0(n5), .B1(n95), .C0(n94), .Y(dout[1])
         );
  AOI2BB2X1 U77 ( .B0(n93), .B1(n112), .A0N(n133), .A1N(n12), .Y(n94) );
  OAI211X1 U78 ( .A0(n128), .A1(n85), .B0(n127), .C0(n126), .Y(dout[3]) );
  AOI32XL U79 ( .A0(n125), .A1(n1), .A2(n124), .B0(n123), .B1(n136), .Y(n126)
         );
  OAI31X1 U80 ( .A0(n122), .A1(n121), .A2(n120), .B0(n85), .Y(n127) );
  OAI221X1 U81 ( .A0(n3), .A1(n108), .B0(n107), .B1(n16), .C0(n106), .Y(
        dout[2]) );
  AOI32XL U82 ( .A0(n105), .A1(n85), .A2(n140), .B0(n2), .B1(n104), .Y(n106)
         );
  AOI211X1 U83 ( .A0(n101), .A1(n4), .B0(n100), .C0(n99), .Y(n107) );
  NAND2X1 U84 ( .A(n148), .B(n147), .Y(dout[4]) );
  AOI222XL U85 ( .A0(n136), .A1(n141), .B0(n3), .B1(n135), .C0(n134), .C1(n138), .Y(n148) );
  AOI222XL U86 ( .A0(n5), .A1(n146), .B0(n145), .B1(n144), .C0(n143), .C1(n85), 
        .Y(n147) );
  CLKINVX3 U87 ( .A(n3), .Y(n16) );
  CLKINVX3 U88 ( .A(n4), .Y(n83) );
  CLKINVX3 U89 ( .A(n5), .Y(n85) );
  CLKINVX3 U90 ( .A(addr[1]), .Y(n86) );
  CLKINVX3 U91 ( .A(addr[3]), .Y(n87) );
endmodule


module sbox8_2 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132;

  NAND2X2 U41 ( .A(addr[6]), .B(n75), .Y(n131) );
  NAND2X2 U48 ( .A(addr[4]), .B(n9), .Y(n123) );
  NAND2X2 U49 ( .A(n2), .B(n12), .Y(n87) );
  NAND2X2 U50 ( .A(addr[1]), .B(n15), .Y(n124) );
  NAND2X2 U54 ( .A(addr[2]), .B(n6), .Y(n116) );
  NAND2X2 U60 ( .A(addr[6]), .B(addr[1]), .Y(n105) );
  NAND2X2 U61 ( .A(n75), .B(n15), .Y(n108) );
  OAI32X1 U1 ( .A0(n15), .A1(addr[4]), .A2(n92), .B0(n115), .B1(n108), .Y(n96)
         );
  OAI31X1 U2 ( .A0(n123), .A1(addr[6]), .A2(n116), .B0(n109), .Y(n110) );
  AOI222X1 U3 ( .A0(n88), .A1(addr[2]), .B0(n12), .B1(n7), .C0(n10), .C1(n92), 
        .Y(n114) );
  OAI222X1 U4 ( .A0(addr[2]), .A1(n126), .B0(n9), .B1(n125), .C0(n124), .C1(
        n123), .Y(n127) );
  OAI221X1 U5 ( .A0(n105), .A1(n87), .B0(addr[4]), .B1(n108), .C0(n86), .Y(n90) );
  NAND2X4 U6 ( .A(addr[4]), .B(n2), .Y(n115) );
  AOI32XL U7 ( .A0(n13), .A1(n5), .A2(n2), .B0(n14), .B1(n117), .Y(n130) );
  OA21XL U8 ( .A0(n10), .A1(n6), .B0(n121), .Y(n78) );
  INVXL U9 ( .A(n119), .Y(n3) );
  INVX3 U10 ( .A(n2), .Y(n9) );
  BUFX4 U11 ( .A(addr[3]), .Y(n2) );
  CLKBUFX3 U12 ( .A(addr[5]), .Y(n1) );
  CLKINVX1 U13 ( .A(n108), .Y(n14) );
  CLKINVX1 U14 ( .A(n107), .Y(n4) );
  CLKINVX1 U15 ( .A(n93), .Y(n8) );
  NAND2X1 U16 ( .A(n9), .B(n12), .Y(n93) );
  NAND2X1 U17 ( .A(n10), .B(n6), .Y(n121) );
  OAI21XL U18 ( .A0(n115), .A1(n6), .B0(n107), .Y(n77) );
  OAI21X1 U19 ( .A0(n12), .A1(n6), .B0(n123), .Y(n88) );
  OAI31XL U20 ( .A0(n115), .A1(n75), .A2(n116), .B0(n118), .Y(n94) );
  CLKINVX1 U21 ( .A(n131), .Y(n74) );
  NAND2X1 U22 ( .A(n5), .B(n9), .Y(n107) );
  OAI22XL U23 ( .A0(n116), .A1(n123), .B0(n5), .B1(n115), .Y(n117) );
  OAI22XL U24 ( .A0(n123), .A1(n108), .B0(n131), .B1(n93), .Y(n95) );
  OAI2BB2XL U25 ( .B0(n115), .B1(n131), .A0N(n88), .A1N(n16), .Y(n89) );
  AOI211XL U26 ( .A0(n108), .A1(n105), .B0(n12), .C0(n121), .Y(n85) );
  CLKINVX1 U27 ( .A(n124), .Y(n13) );
  OAI22XL U28 ( .A0(n5), .A1(n123), .B0(n78), .B1(n87), .Y(n81) );
  NAND2BX2 U29 ( .AN(n78), .B(n9), .Y(n120) );
  NAND2XL U30 ( .A(n115), .B(n93), .Y(n104) );
  OAI2BB2XL U31 ( .B0(n106), .B1(n105), .A0N(n104), .A1N(n13), .Y(n111) );
  NOR2BXL U32 ( .AN(n123), .B(n103), .Y(n106) );
  NAND3X1 U33 ( .A(n104), .B(n75), .C(n5), .Y(n84) );
  AO21X1 U34 ( .A0(n5), .A1(n16), .B0(n101), .Y(n102) );
  OAI33X1 U35 ( .A0(n15), .A1(n9), .A2(n100), .B0(n10), .B1(n103), .B2(n124), 
        .Y(n101) );
  OA22XL U36 ( .A0(n107), .A1(n131), .B0(n120), .B1(n124), .Y(n98) );
  CLKINVX1 U37 ( .A(n125), .Y(n11) );
  OAI21XL U38 ( .A0(n13), .A1(n74), .B0(addr[4]), .Y(n86) );
  NAND2X1 U39 ( .A(n1), .B(n10), .Y(n100) );
  OAI221X1 U40 ( .A0(n124), .A1(n121), .B0(addr[1]), .B1(n120), .C0(n3), .Y(
        n128) );
  OAI31XL U42 ( .A0(n10), .A1(n75), .A2(n9), .B0(n118), .Y(n119) );
  NAND2X1 U43 ( .A(n16), .B(addr[2]), .Y(n125) );
  NAND4XL U44 ( .A(n74), .B(n1), .C(n2), .D(addr[2]), .Y(n109) );
  NAND3X1 U45 ( .A(n5), .B(n15), .C(n2), .Y(n118) );
  OAI21XL U46 ( .A0(n1), .A1(n87), .B0(n114), .Y(n76) );
  OAI22XL U47 ( .A0(n108), .A1(n120), .B0(n79), .B1(n100), .Y(n80) );
  AOI221XL U51 ( .A0(n74), .A1(n9), .B0(n16), .B1(n2), .C0(n91), .Y(n79) );
  NOR2X1 U52 ( .A(n1), .B(n2), .Y(n103) );
  NOR2X1 U53 ( .A(n87), .B(addr[6]), .Y(n91) );
  NOR2X1 U55 ( .A(n9), .B(n1), .Y(n92) );
  CLKINVX1 U56 ( .A(n100), .Y(n7) );
  OA21XL U57 ( .A0(n1), .A1(n115), .B0(n120), .Y(n132) );
  AOI221XL U58 ( .A0(n14), .A1(n2), .B0(n16), .B1(addr[4]), .C0(n122), .Y(n126) );
  OAI22XL U59 ( .A0(n2), .A1(n75), .B0(addr[4]), .B1(n131), .Y(n122) );
  OAI211X1 U62 ( .A0(addr[2]), .A1(n99), .B0(n98), .C0(n97), .Y(dout[2]) );
  AOI221XL U63 ( .A0(addr[2]), .A1(n96), .B0(n1), .B1(n95), .C0(n94), .Y(n97)
         );
  AOI221XL U64 ( .A0(n91), .A1(n1), .B0(n90), .B1(n6), .C0(n89), .Y(n99) );
  OAI211X1 U65 ( .A0(n132), .A1(n131), .B0(n130), .C0(n129), .Y(dout[4]) );
  AOI222XL U66 ( .A0(n128), .A1(n12), .B0(n1), .B1(n127), .C0(n4), .C1(n16), 
        .Y(n129) );
  OAI211X1 U67 ( .A0(addr[1]), .A1(n114), .B0(n113), .C0(n112), .Y(dout[3]) );
  AOI221XL U68 ( .A0(n111), .A1(n10), .B0(n4), .B1(n14), .C0(n110), .Y(n112)
         );
  AOI2BB2XL U69 ( .B0(n102), .B1(n12), .A0N(n115), .A1N(n125), .Y(n113) );
  NAND4BX1 U70 ( .AN(n85), .B(n84), .C(n83), .D(n82), .Y(dout[1]) );
  AOI221XL U71 ( .A0(n74), .A1(n81), .B0(n8), .B1(n11), .C0(n80), .Y(n82) );
  AOI22X1 U72 ( .A0(n16), .A1(n77), .B0(n13), .B1(n76), .Y(n83) );
  CLKINVX3 U73 ( .A(n116), .Y(n5) );
  CLKINVX3 U74 ( .A(n1), .Y(n6) );
  CLKINVX3 U75 ( .A(addr[2]), .Y(n10) );
  CLKINVX3 U76 ( .A(addr[4]), .Y(n12) );
  CLKINVX3 U77 ( .A(addr[6]), .Y(n15) );
  CLKINVX3 U78 ( .A(n105), .Y(n16) );
  CLKINVX3 U79 ( .A(addr[1]), .Y(n75) );
endmodule


module crp_2 ( P, R, K_sub );
  output [1:32] P;
  input [1:32] R;
  input [1:48] K_sub;
  wire   n1;
  wire   [1:48] X;

  sbox1_2 u0 ( .addr(X[1:6]), .dout({P[9], P[17], P[23], P[31]}) );
  sbox2_2 u1 ( .addr({X[7], n1, X[9:12]}), .dout({P[13], P[28], P[2], P[18]})
         );
  sbox3_2 u2 ( .addr(X[13:18]), .dout({P[24], P[16], P[30], P[6]}) );
  sbox4_2 u3 ( .addr(X[19:24]), .dout({P[26], P[20], P[10], P[1]}) );
  sbox5_2 u4 ( .addr(X[25:30]), .dout({P[8], P[14], P[25], P[3]}) );
  sbox6_2 u5 ( .addr(X[31:36]), .dout({P[4], P[29], P[11], P[19]}) );
  sbox7_2 u6 ( .addr(X[37:42]), .dout({P[32], P[12], P[22], P[7]}) );
  sbox8_2 u7 ( .addr(X[43:48]), .dout({P[5], P[27], P[15], P[21]}) );
  XNOR2X1 U1 ( .A(R[5]), .B(K_sub[8]), .Y(X[8]) );
  INVX3 U2 ( .A(X[8]), .Y(n1) );
  XOR2X1 U3 ( .A(R[1]), .B(K_sub[2]), .Y(X[2]) );
  CLKXOR2X4 U4 ( .A(R[29]), .B(K_sub[42]), .Y(X[42]) );
  CLKXOR2X4 U5 ( .A(R[16]), .B(K_sub[25]), .Y(X[25]) );
  CLKXOR2X4 U6 ( .A(R[8]), .B(K_sub[11]), .Y(X[11]) );
  CLKXOR2X4 U7 ( .A(R[22]), .B(K_sub[33]), .Y(X[33]) );
  CLKXOR2X4 U8 ( .A(R[29]), .B(K_sub[44]), .Y(X[44]) );
  CLKXOR2X4 U9 ( .A(R[16]), .B(K_sub[23]), .Y(X[23]) );
  CLKXOR2X4 U10 ( .A(R[10]), .B(K_sub[15]), .Y(X[15]) );
  CLKXOR2X4 U11 ( .A(R[20]), .B(K_sub[31]), .Y(X[31]) );
  CLKXOR2X4 U12 ( .A(R[31]), .B(K_sub[46]), .Y(X[46]) );
  CLKXOR2X4 U13 ( .A(R[12]), .B(K_sub[19]), .Y(X[19]) );
  CLKXOR2X4 U14 ( .A(R[26]), .B(K_sub[39]), .Y(X[39]) );
  CLKXOR2X4 U15 ( .A(R[20]), .B(K_sub[29]), .Y(X[29]) );
  CLKXOR2X2 U16 ( .A(R[4]), .B(K_sub[5]), .Y(X[5]) );
  CLKXOR2X2 U17 ( .A(R[15]), .B(K_sub[22]), .Y(X[22]) );
  CLKXOR2X2 U18 ( .A(R[24]), .B(K_sub[35]), .Y(X[35]) );
  CLKXOR2X2 U19 ( .A(R[21]), .B(K_sub[30]), .Y(X[30]) );
  CLKXOR2X2 U20 ( .A(R[12]), .B(K_sub[17]), .Y(X[17]) );
  CLKXOR2X2 U21 ( .A(R[32]), .B(K_sub[1]), .Y(X[1]) );
  CLKXOR2X2 U22 ( .A(R[13]), .B(K_sub[20]), .Y(X[20]) );
  CLKXOR2X2 U23 ( .A(R[18]), .B(K_sub[27]), .Y(X[27]) );
  CLKXOR2X2 U24 ( .A(R[8]), .B(K_sub[13]), .Y(X[13]) );
  CLKXOR2X2 U25 ( .A(R[5]), .B(K_sub[6]), .Y(X[6]) );
  CLKXOR2X2 U26 ( .A(R[4]), .B(K_sub[7]), .Y(X[7]) );
  CLKXOR2X2 U27 ( .A(R[24]), .B(K_sub[37]), .Y(X[37]) );
  CLKXOR2X2 U28 ( .A(R[28]), .B(K_sub[43]), .Y(X[43]) );
  CLKXOR2X2 U29 ( .A(R[1]), .B(K_sub[48]), .Y(X[48]) );
  CLKXOR2X2 U30 ( .A(R[17]), .B(K_sub[24]), .Y(X[24]) );
  CLKXOR2X2 U31 ( .A(R[9]), .B(K_sub[12]), .Y(X[12]) );
  CLKXOR2X2 U32 ( .A(R[13]), .B(K_sub[18]), .Y(X[18]) );
  CLKXOR2X2 U33 ( .A(R[25]), .B(K_sub[36]), .Y(X[36]) );
  XOR2X1 U34 ( .A(R[23]), .B(K_sub[34]), .Y(X[34]) );
  XOR2X1 U35 ( .A(R[9]), .B(K_sub[14]), .Y(X[14]) );
  XOR2X1 U36 ( .A(R[30]), .B(K_sub[45]), .Y(X[45]) );
  XOR2X1 U37 ( .A(R[21]), .B(K_sub[32]), .Y(X[32]) );
  XOR2X1 U38 ( .A(R[25]), .B(K_sub[38]), .Y(X[38]) );
  XOR2X1 U39 ( .A(R[27]), .B(K_sub[40]), .Y(X[40]) );
  XOR2X1 U40 ( .A(R[3]), .B(K_sub[4]), .Y(X[4]) );
  XOR2X1 U41 ( .A(R[11]), .B(K_sub[16]), .Y(X[16]) );
  XOR2X1 U42 ( .A(R[7]), .B(K_sub[10]), .Y(X[10]) );
  XOR2X1 U43 ( .A(R[14]), .B(K_sub[21]), .Y(X[21]) );
  XOR2X1 U44 ( .A(R[6]), .B(K_sub[9]), .Y(X[9]) );
  XOR2X1 U45 ( .A(R[2]), .B(K_sub[3]), .Y(X[3]) );
  XOR2X1 U46 ( .A(R[28]), .B(K_sub[41]), .Y(X[41]) );
  XOR2X1 U47 ( .A(R[17]), .B(K_sub[26]), .Y(X[26]) );
  XOR2X1 U48 ( .A(R[32]), .B(K_sub[47]), .Y(X[47]) );
  XOR2X1 U49 ( .A(R[19]), .B(K_sub[28]), .Y(X[28]) );
endmodule


module sbox1_1 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127;

  OAI222X4 U13 ( .A0(addr[5]), .A1(n101), .B0(n1), .B1(n100), .C0(n99), .C1(
        n72), .Y(dout[3]) );
  OAI21X2 U42 ( .A0(n4), .A1(n112), .B0(n106), .Y(n123) );
  NAND2X2 U44 ( .A(addr[6]), .B(n9), .Y(n115) );
  NAND2X2 U48 ( .A(addr[1]), .B(n12), .Y(n114) );
  OAI22X2 U49 ( .A0(n6), .A1(n71), .B0(addr[5]), .B1(n120), .Y(n85) );
  NAND2X2 U50 ( .A(n3), .B(n6), .Y(n120) );
  NOR2X2 U51 ( .A(n6), .B(n3), .Y(n124) );
  NOR3X2 U55 ( .A(n2), .B(addr[6]), .C(n72), .Y(n102) );
  NOR2X2 U56 ( .A(n109), .B(n3), .Y(n93) );
  NAND2X2 U57 ( .A(addr[1]), .B(addr[6]), .Y(n109) );
  NAND2X2 U59 ( .A(n9), .B(n12), .Y(n112) );
  NOR2X1 U1 ( .A(n114), .B(n120), .Y(n104) );
  BUFX4 U2 ( .A(addr[4]), .Y(n2) );
  CLKBUFX3 U3 ( .A(addr[2]), .Y(n1) );
  OAI32X1 U4 ( .A0(n112), .A1(n2), .A2(n4), .B0(n115), .B1(n113), .Y(n80) );
  NOR2BXL U5 ( .AN(n118), .B(n1), .Y(n122) );
  CLKBUFX3 U6 ( .A(addr[2]), .Y(n4) );
  INVX3 U7 ( .A(addr[6]), .Y(n12) );
  OAI221X4 U8 ( .A0(n88), .A1(n71), .B0(addr[5]), .B1(n87), .C0(n86), .Y(
        dout[2]) );
  OAI221X4 U9 ( .A0(addr[5]), .A1(n127), .B0(n126), .B1(n71), .C0(n125), .Y(
        dout[4]) );
  OA21XL U10 ( .A0(n95), .A1(n115), .B0(n107), .Y(n119) );
  AOI222XL U11 ( .A0(n8), .A1(n1), .B0(n2), .B1(n110), .C0(n10), .C1(n72), .Y(
        n111) );
  AOI2BB2X1 U12 ( .B0(n2), .B1(n10), .A0N(addr[4]), .A1N(n115), .Y(n91) );
  BUFX4 U14 ( .A(addr[3]), .Y(n3) );
  CLKINVX1 U15 ( .A(n112), .Y(n8) );
  CLKINVX1 U16 ( .A(n113), .Y(n13) );
  NAND2BX1 U17 ( .AN(n104), .B(n119), .Y(n84) );
  CLKXOR2X2 U18 ( .A(n69), .B(n72), .Y(n90) );
  NOR2X1 U19 ( .A(n6), .B(n69), .Y(n118) );
  OAI21XL U20 ( .A0(n69), .A1(n114), .B0(n91), .Y(n92) );
  NAND2X1 U21 ( .A(n93), .B(n6), .Y(n107) );
  NAND2X1 U22 ( .A(n72), .B(n69), .Y(n113) );
  OAI211X1 U23 ( .A0(n6), .A1(n114), .B0(n108), .C0(n107), .Y(n89) );
  CLKINVX1 U24 ( .A(n109), .Y(n10) );
  NAND2X1 U25 ( .A(n124), .B(n7), .Y(n108) );
  CLKINVX1 U26 ( .A(n114), .Y(n11) );
  CLKINVX1 U27 ( .A(n115), .Y(n7) );
  CLKINVX1 U28 ( .A(n95), .Y(n70) );
  AO22X1 U29 ( .A0(n90), .A1(n7), .B0(n69), .B1(n123), .Y(n76) );
  OAI31X1 U30 ( .A0(n72), .A1(n3), .A2(n9), .B0(n103), .Y(n105) );
  AOI31XL U31 ( .A0(n9), .A1(n72), .A2(n2), .B0(n102), .Y(n103) );
  AOI211X1 U32 ( .A0(n5), .A1(n4), .B0(n117), .C0(n116), .Y(n126) );
  CLKINVX1 U33 ( .A(n108), .Y(n5) );
  AOI211X1 U34 ( .A0(n115), .A1(n114), .B0(n113), .C0(n2), .Y(n116) );
  OAI22X1 U35 ( .A0(n120), .A1(n112), .B0(n111), .B1(n69), .Y(n117) );
  AOI211X1 U36 ( .A0(n10), .A1(n118), .B0(n81), .C0(n80), .Y(n88) );
  OAI22X1 U37 ( .A0(n91), .A1(n72), .B0(n3), .B1(n106), .Y(n81) );
  CLKINVX3 U38 ( .A(addr[5]), .Y(n71) );
  NAND2X1 U39 ( .A(n3), .B(n71), .Y(n95) );
  NAND2X1 U40 ( .A(n11), .B(n1), .Y(n106) );
  XOR2X1 U41 ( .A(n82), .B(n2), .Y(n83) );
  NAND2X1 U43 ( .A(n1), .B(n3), .Y(n82) );
  OAI22XL U45 ( .A0(n3), .A1(n9), .B0(n69), .B1(n112), .Y(n94) );
  AOI211XL U46 ( .A0(n98), .A1(n69), .B0(n97), .C0(n104), .Y(n99) );
  OAI22XL U47 ( .A0(n96), .A1(n6), .B0(n95), .B1(n109), .Y(n97) );
  OAI22XL U52 ( .A0(n12), .A1(n71), .B0(n2), .B1(addr[1]), .Y(n98) );
  AOI221XL U53 ( .A0(n70), .A1(addr[6]), .B0(addr[5]), .B1(n94), .C0(n93), .Y(
        n96) );
  OAI21XL U54 ( .A0(addr[1]), .A1(n120), .B0(n119), .Y(n121) );
  AOI221XL U58 ( .A0(n8), .A1(n118), .B0(n93), .B1(n71), .C0(n75), .Y(n78) );
  OAI31X1 U60 ( .A0(n71), .A1(n2), .A2(n74), .B0(n73), .Y(n75) );
  OA21XL U61 ( .A0(n3), .A1(n12), .B0(n109), .Y(n74) );
  OAI21XL U62 ( .A0(n124), .A1(n85), .B0(n11), .Y(n73) );
  OAI21XL U63 ( .A0(n1), .A1(n9), .B0(n109), .Y(n110) );
  INVX4 U64 ( .A(n4), .Y(n72) );
  AOI32X1 U65 ( .A0(n4), .A1(n85), .A2(n8), .B0(n84), .B1(n72), .Y(n86) );
  AOI222XL U66 ( .A0(n124), .A1(n9), .B0(n83), .B1(addr[1]), .C0(n13), .C1(n12), .Y(n87) );
  OAI221X1 U67 ( .A0(n79), .A1(n71), .B0(n4), .B1(n78), .C0(n77), .Y(dout[1])
         );
  AOI32XL U68 ( .A0(addr[6]), .A1(n85), .A2(n1), .B0(n76), .B1(n71), .Y(n77)
         );
  AOI221X1 U69 ( .A0(n8), .A1(n90), .B0(n4), .B1(n93), .C0(n102), .Y(n79) );
  AOI222XL U70 ( .A0(n124), .A1(n123), .B0(n122), .B1(addr[6]), .C0(n1), .C1(
        n121), .Y(n125) );
  NOR4BBX1 U71 ( .AN(n107), .BN(n106), .C(n105), .D(n104), .Y(n127) );
  AOI222XL U72 ( .A0(n8), .A1(n90), .B0(n89), .B1(n72), .C0(n123), .C1(n6), 
        .Y(n101) );
  AOI2BB2XL U73 ( .B0(addr[5]), .B1(n92), .A0N(n120), .A1N(addr[1]), .Y(n100)
         );
  CLKINVX3 U74 ( .A(n2), .Y(n6) );
  CLKINVX3 U75 ( .A(addr[1]), .Y(n9) );
  CLKINVX3 U76 ( .A(n3), .Y(n69) );
endmodule


module sbox2_1 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147;

  NAND2X2 U55 ( .A(n2), .B(n6), .Y(n136) );
  NAND2X2 U57 ( .A(addr[2]), .B(n11), .Y(n104) );
  NAND2X2 U60 ( .A(addr[5]), .B(addr[2]), .Y(n132) );
  NOR2X2 U61 ( .A(n16), .B(n13), .Y(n101) );
  NAND2X2 U62 ( .A(n15), .B(n83), .Y(n146) );
  NAND2X2 U63 ( .A(n3), .B(n82), .Y(n124) );
  NAND2X2 U64 ( .A(addr[6]), .B(n15), .Y(n122) );
  NAND2X2 U67 ( .A(n3), .B(n2), .Y(n133) );
  CLKINVX1 U1 ( .A(n121), .Y(n16) );
  AOI222XL U2 ( .A0(n5), .A1(n81), .B0(n88), .B1(n82), .C0(n140), .C1(n13), 
        .Y(n89) );
  AOI211X1 U3 ( .A0(n12), .A1(n95), .B0(n94), .C0(n93), .Y(n96) );
  CLKINVX1 U4 ( .A(addr[5]), .Y(n1) );
  OAI22X1 U5 ( .A0(n117), .A1(n114), .B0(n89), .B1(n11), .Y(n94) );
  INVX3 U6 ( .A(addr[5]), .Y(n11) );
  OAI211X4 U7 ( .A0(n147), .A1(n146), .B0(n145), .C0(n144), .Y(dout[4]) );
  NAND2X1 U8 ( .A(addr[1]), .B(addr[6]), .Y(n121) );
  CLKINVX2 U9 ( .A(addr[1]), .Y(n15) );
  OAI221X1 U10 ( .A0(addr[1]), .A1(n136), .B0(n133), .B1(n15), .C0(n87), .Y(
        n95) );
  NOR2X1 U11 ( .A(n104), .B(n2), .Y(n141) );
  NOR2X1 U12 ( .A(n124), .B(n2), .Y(n140) );
  CLKBUFX4 U13 ( .A(addr[4]), .Y(n2) );
  NAND2X4 U14 ( .A(addr[1]), .B(n83), .Y(n114) );
  INVX3 U15 ( .A(addr[6]), .Y(n83) );
  NAND2XL U16 ( .A(n102), .B(n6), .Y(n109) );
  AOI2BB2X1 U17 ( .B0(n11), .B1(n8), .A0N(n104), .A1N(n136), .Y(n117) );
  NOR3BXL U18 ( .AN(n135), .B(n134), .C(n5), .Y(n147) );
  BUFX4 U19 ( .A(addr[3]), .Y(n3) );
  NAND2X1 U20 ( .A(n5), .B(n16), .Y(n113) );
  CLKINVX1 U21 ( .A(n146), .Y(n13) );
  CLKINVX1 U22 ( .A(n115), .Y(n5) );
  CLKINVX1 U23 ( .A(n122), .Y(n14) );
  OAI31X1 U24 ( .A0(n124), .A1(n83), .A2(n11), .B0(n123), .Y(n128) );
  OAI21XL U25 ( .A0(n1), .A1(n15), .B0(n140), .Y(n123) );
  OAI22X1 U26 ( .A0(n122), .A1(n124), .B0(n101), .B1(n132), .Y(n84) );
  INVX1 U27 ( .A(n114), .Y(n81) );
  OAI22X1 U28 ( .A0(n122), .A1(n6), .B0(n9), .B1(n121), .Y(n129) );
  NAND3X1 U29 ( .A(n9), .B(n11), .C(n15), .Y(n111) );
  NAND2X1 U30 ( .A(n6), .B(n9), .Y(n115) );
  OAI21XL U31 ( .A0(n82), .A1(n133), .B0(n135), .Y(n85) );
  OAI22XL U32 ( .A0(n117), .A1(n146), .B0(n116), .B1(n132), .Y(n118) );
  AOI222XL U33 ( .A0(n81), .A1(n115), .B0(n7), .B1(n83), .C0(n5), .C1(n13), 
        .Y(n116) );
  CLKINVX1 U34 ( .A(n104), .Y(n10) );
  OAI2BB2XL U35 ( .B0(n114), .B1(n135), .A0N(n126), .A1N(n7), .Y(n106) );
  OAI21XL U36 ( .A0(n112), .A1(n114), .B0(n111), .Y(n120) );
  OAI21XL U37 ( .A0(n133), .A1(n114), .B0(n113), .Y(n119) );
  CLKINVX1 U38 ( .A(n124), .Y(n8) );
  CLKINVX1 U39 ( .A(n136), .Y(n4) );
  CLKINVX1 U40 ( .A(n133), .Y(n7) );
  CLKINVX1 U41 ( .A(n132), .Y(n12) );
  AOI2BB1X1 U42 ( .A0N(n126), .A1N(n125), .B0(n136), .Y(n127) );
  OAI22XL U43 ( .A0(n104), .A1(n114), .B0(n101), .B1(n132), .Y(n102) );
  AO21XL U44 ( .A0(n82), .A1(n4), .B0(n141), .Y(n86) );
  AO21X1 U45 ( .A0(n6), .A1(n10), .B0(n140), .Y(n142) );
  NAND3X1 U46 ( .A(n82), .B(n9), .C(addr[5]), .Y(n135) );
  OAI22X1 U47 ( .A0(addr[5]), .A1(n121), .B0(n122), .B1(n11), .Y(n126) );
  AOI2BB1X1 U48 ( .A0N(n3), .A1N(n1), .B0(n4), .Y(n112) );
  NOR3X1 U49 ( .A(addr[1]), .B(addr[2]), .C(n11), .Y(n125) );
  AOI2BB1XL U50 ( .A0N(n92), .A1N(n91), .B0(addr[5]), .Y(n93) );
  OAI31XL U51 ( .A0(n114), .A1(n2), .A2(n6), .B0(n90), .Y(n91) );
  OAI21XL U52 ( .A0(n7), .A1(n8), .B0(n14), .Y(n90) );
  NAND2X1 U53 ( .A(n81), .B(n2), .Y(n137) );
  OAI31XL U54 ( .A0(n101), .A1(n3), .A2(addr[2]), .B0(n113), .Y(n92) );
  OAI211X1 U56 ( .A0(n139), .A1(n11), .B0(n138), .C0(n137), .Y(n143) );
  NAND3X1 U58 ( .A(n9), .B(n11), .C(addr[6]), .Y(n138) );
  AOI2BB2X1 U59 ( .B0(n14), .B1(n6), .A0N(n15), .A1N(n136), .Y(n139) );
  OAI22XL U65 ( .A0(addr[5]), .A1(n133), .B0(n3), .B1(n132), .Y(n134) );
  OAI2BB2XL U66 ( .B0(n112), .B1(n122), .A0N(n1), .A1N(n99), .Y(n100) );
  OAI211X1 U68 ( .A0(n146), .A1(n2), .B0(n137), .C0(n113), .Y(n99) );
  NAND3X1 U69 ( .A(n14), .B(n9), .C(n3), .Y(n87) );
  AOI2BB2XL U70 ( .B0(n3), .B1(n105), .A0N(n137), .A1N(n132), .Y(n108) );
  OAI211XL U71 ( .A0(n104), .A1(n146), .B0(n103), .C0(n111), .Y(n105) );
  NAND3XL U72 ( .A(addr[5]), .B(n9), .C(n16), .Y(n103) );
  OAI22XL U73 ( .A0(n3), .A1(n114), .B0(n83), .B1(n115), .Y(n88) );
  AOI33XL U74 ( .A0(n14), .A1(n10), .A2(n2), .B0(n12), .B1(n146), .B2(n3), .Y(
        n145) );
  AOI222XL U75 ( .A0(n143), .A1(n82), .B0(n16), .B1(n142), .C0(n81), .C1(n141), 
        .Y(n144) );
  NAND2X1 U76 ( .A(n131), .B(n130), .Y(dout[3]) );
  AOI221XL U77 ( .A0(n120), .A1(n82), .B0(addr[2]), .B1(n119), .C0(n118), .Y(
        n131) );
  AOI211X1 U78 ( .A0(n10), .A1(n129), .B0(n128), .C0(n127), .Y(n130) );
  NAND4X1 U79 ( .A(n110), .B(n109), .C(n108), .D(n107), .Y(dout[2]) );
  AOI32XL U80 ( .A0(addr[1]), .A1(addr[2]), .A2(n4), .B0(n100), .B1(n82), .Y(
        n110) );
  AOI221XL U81 ( .A0(n125), .A1(addr[4]), .B0(n141), .B1(n14), .C0(n106), .Y(
        n107) );
  NAND3X1 U82 ( .A(n98), .B(n97), .C(n96), .Y(dout[1]) );
  AOI32XL U83 ( .A0(n10), .A1(n15), .A2(n5), .B0(n13), .B1(n86), .Y(n97) );
  AOI22X1 U84 ( .A0(n16), .A1(n85), .B0(n2), .B1(n84), .Y(n98) );
  CLKINVX3 U85 ( .A(n3), .Y(n6) );
  CLKINVX3 U86 ( .A(n2), .Y(n9) );
  CLKINVX3 U87 ( .A(addr[2]), .Y(n82) );
endmodule


module sbox3_1 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134;

  NOR2X2 U35 ( .A(n17), .B(addr[3]), .Y(n109) );
  NOR2X2 U50 ( .A(addr[1]), .B(addr[6]), .Y(n108) );
  NOR2X2 U52 ( .A(n77), .B(n3), .Y(n88) );
  NOR2X2 U56 ( .A(n77), .B(n78), .Y(n95) );
  NOR2X1 U1 ( .A(n17), .B(n77), .Y(n107) );
  OAI221X1 U2 ( .A0(n125), .A1(n17), .B0(n4), .B1(addr[1]), .C0(n14), .Y(n105)
         );
  INVXL U3 ( .A(n2), .Y(n1) );
  NOR2X1 U4 ( .A(n10), .B(n4), .Y(n92) );
  NOR2X1 U5 ( .A(n19), .B(n4), .Y(n122) );
  NOR2X1 U6 ( .A(n14), .B(n4), .Y(n96) );
  CLKBUFX3 U7 ( .A(addr[2]), .Y(n4) );
  INVX1 U8 ( .A(addr[2]), .Y(n2) );
  NOR2X1 U9 ( .A(n4), .B(n3), .Y(n111) );
  BUFX4 U10 ( .A(addr[4]), .Y(n3) );
  OAI33X1 U11 ( .A0(n19), .A1(n126), .A2(n78), .B0(n17), .B1(n95), .B2(n120), 
        .Y(n80) );
  INVX3 U12 ( .A(n4), .Y(n78) );
  OAI221X1 U13 ( .A0(addr[5]), .A1(n91), .B0(n90), .B1(n79), .C0(n89), .Y(
        dout[1]) );
  NOR2X4 U14 ( .A(n11), .B(n15), .Y(n125) );
  NOR2X4 U15 ( .A(addr[3]), .B(n3), .Y(n131) );
  NOR2X4 U16 ( .A(n15), .B(addr[6]), .Y(n126) );
  INVX3 U17 ( .A(addr[1]), .Y(n15) );
  NAND2XL U18 ( .A(n95), .B(n125), .Y(n133) );
  OAI211XL U19 ( .A0(n3), .A1(n9), .B0(n129), .C0(n128), .Y(n130) );
  NAND4XL U20 ( .A(n115), .B(n114), .C(n113), .D(n112), .Y(n116) );
  CLKINVX1 U21 ( .A(n133), .Y(n7) );
  INVX1 U22 ( .A(n125), .Y(n5) );
  CLKINVX1 U23 ( .A(n107), .Y(n16) );
  NAND2X1 U24 ( .A(n10), .B(n12), .Y(n123) );
  CLKINVX1 U25 ( .A(n87), .Y(n12) );
  CLKINVX1 U26 ( .A(n121), .Y(n76) );
  CLKINVX1 U27 ( .A(n120), .Y(n6) );
  CLKINVX1 U28 ( .A(n115), .Y(n8) );
  CLKINVX1 U29 ( .A(n108), .Y(n14) );
  NOR2X1 U30 ( .A(n10), .B(n78), .Y(n104) );
  NOR2X1 U31 ( .A(n5), .B(n78), .Y(n110) );
  INVX1 U32 ( .A(n126), .Y(n13) );
  AOI21X1 U33 ( .A0(n77), .A1(n78), .B0(n95), .Y(n121) );
  OAI21XL U34 ( .A0(n111), .A1(n131), .B0(n125), .Y(n83) );
  CLKINVX1 U36 ( .A(n82), .Y(n10) );
  NOR2X1 U37 ( .A(n13), .B(n17), .Y(n87) );
  NOR2X1 U38 ( .A(n125), .B(n108), .Y(n120) );
  OAI21XL U39 ( .A0(n110), .A1(n92), .B0(n131), .Y(n101) );
  NAND2X1 U40 ( .A(n104), .B(n88), .Y(n115) );
  CLKINVX1 U41 ( .A(n88), .Y(n19) );
  CLKINVX1 U42 ( .A(n92), .Y(n9) );
  CLKINVX1 U43 ( .A(n111), .Y(n20) );
  CLKINVX1 U44 ( .A(n122), .Y(n18) );
  OR2X1 U45 ( .A(n104), .B(n96), .Y(n127) );
  OAI221X1 U46 ( .A0(n13), .A1(n20), .B0(n78), .B1(n12), .C0(n94), .Y(n99) );
  AOI221XL U47 ( .A0(n96), .A1(n3), .B0(n93), .B1(n17), .C0(n7), .Y(n94) );
  OAI21XL U48 ( .A0(n78), .A1(n14), .B0(n9), .Y(n93) );
  XNOR2X1 U49 ( .A(addr[5]), .B(addr[3]), .Y(n103) );
  CLKINVX1 U51 ( .A(addr[5]), .Y(n79) );
  OAI221X1 U53 ( .A0(n14), .A1(n20), .B0(n5), .B1(n19), .C0(n106), .Y(n117) );
  AOI221XL U54 ( .A0(addr[3]), .A1(n105), .B0(n104), .B1(n131), .C0(n7), .Y(
        n106) );
  CLKINVX1 U55 ( .A(addr[6]), .Y(n11) );
  NAND3X1 U57 ( .A(n4), .B(n15), .C(n109), .Y(n114) );
  NOR2X1 U58 ( .A(n11), .B(addr[1]), .Y(n82) );
  AOI32XL U59 ( .A0(n78), .A1(n77), .A2(n125), .B0(n124), .B1(n11), .Y(n129)
         );
  AOI22XL U60 ( .A0(n3), .A1(n127), .B0(n126), .B1(n131), .Y(n128) );
  OAI22XL U61 ( .A0(n3), .A1(n2), .B0(n4), .B1(n16), .Y(n124) );
  AOI222XL U62 ( .A0(n111), .A1(n126), .B0(n110), .B1(n77), .C0(n109), .C1(
        n108), .Y(n112) );
  OAI211XL U63 ( .A0(n107), .A1(n131), .B0(n2), .C0(addr[6]), .Y(n113) );
  OAI21XL U64 ( .A0(n1), .A1(addr[1]), .B0(n13), .Y(n81) );
  AOI221XL U65 ( .A0(n87), .A1(n77), .B0(n88), .B1(n126), .C0(n86), .Y(n90) );
  OAI211X1 U66 ( .A0(n85), .A1(n78), .B0(n84), .C0(n83), .Y(n86) );
  AOI222XL U67 ( .A0(n82), .A1(n77), .B0(n108), .B1(n107), .C0(n131), .C1(n15), 
        .Y(n85) );
  OAI21XL U68 ( .A0(n92), .A1(n7), .B0(addr[4]), .Y(n84) );
  AOI221XL U69 ( .A0(n126), .A1(n76), .B0(addr[3]), .B1(n127), .C0(n97), .Y(
        n98) );
  OAI22X1 U70 ( .A0(n5), .A1(n18), .B0(n16), .B1(n10), .Y(n97) );
  OAI211X1 U71 ( .A0(n14), .A1(n18), .B0(n119), .C0(n118), .Y(dout[3]) );
  AOI32XL U72 ( .A0(n126), .A1(n4), .A2(n103), .B0(n109), .B1(n110), .Y(n119)
         );
  AOI22XL U73 ( .A0(n117), .A1(n79), .B0(addr[5]), .B1(n116), .Y(n118) );
  OAI221X1 U74 ( .A0(n134), .A1(n79), .B0(n3), .B1(n133), .C0(n132), .Y(
        dout[4]) );
  AOI32XL U75 ( .A0(n131), .A1(n11), .A2(n1), .B0(n130), .B1(n79), .Y(n132) );
  AOI222XL U76 ( .A0(n76), .A1(n123), .B0(n122), .B1(addr[1]), .C0(n121), .C1(
        n6), .Y(n134) );
  AOI221XL U77 ( .A0(n122), .A1(n126), .B0(n96), .B1(n109), .C0(n8), .Y(n89)
         );
  AOI221XL U78 ( .A0(n131), .A1(n81), .B0(n95), .B1(n123), .C0(n80), .Y(n91)
         );
  NAND4X1 U79 ( .A(n102), .B(n114), .C(n101), .D(n100), .Y(dout[2]) );
  NAND3XL U80 ( .A(n3), .B(n125), .C(n103), .Y(n102) );
  AOI2BB2XL U81 ( .B0(addr[5]), .B1(n99), .A0N(addr[5]), .A1N(n98), .Y(n100)
         );
  CLKINVX3 U82 ( .A(n3), .Y(n17) );
  CLKINVX3 U83 ( .A(addr[3]), .Y(n77) );
endmodule


module sbox4_1 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126;

  OAI32X4 U12 ( .A0(n13), .A1(n2), .A2(addr[2]), .B0(n12), .B1(n108), .Y(n123)
         );
  OAI222X4 U20 ( .A0(addr[2]), .A1(n92), .B0(n106), .B1(n91), .C0(n90), .C1(n4), .Y(dout[2]) );
  OAI222X4 U33 ( .A0(addr[4]), .A1(n106), .B0(n7), .B1(n108), .C0(n2), .C1(
        n118), .Y(n83) );
  NAND2X2 U34 ( .A(addr[4]), .B(n2), .Y(n108) );
  NOR2X2 U43 ( .A(n71), .B(addr[4]), .Y(n113) );
  NOR2X2 U45 ( .A(n12), .B(n2), .Y(n111) );
  NAND2X2 U51 ( .A(n7), .B(n72), .Y(n118) );
  NOR2X2 U52 ( .A(n16), .B(addr[5]), .Y(n97) );
  NAND2X2 U53 ( .A(addr[6]), .B(addr[1]), .Y(n85) );
  NAND2X2 U54 ( .A(addr[1]), .B(n72), .Y(n116) );
  NOR2X2 U55 ( .A(n115), .B(n12), .Y(n121) );
  NAND2X2 U56 ( .A(n71), .B(n16), .Y(n115) );
  NAND2X2 U57 ( .A(addr[5]), .B(n16), .Y(n96) );
  NAND2X2 U58 ( .A(addr[6]), .B(n7), .Y(n106) );
  OAI222X1 U1 ( .A0(n13), .A1(n85), .B0(n97), .B1(n116), .C0(n16), .C1(n118), 
        .Y(n73) );
  CLKINVX1 U2 ( .A(n116), .Y(n10) );
  CLKINVX1 U3 ( .A(n71), .Y(n1) );
  CLKBUFX3 U4 ( .A(addr[3]), .Y(n2) );
  OAI31X4 U5 ( .A0(n118), .A1(n12), .A2(n16), .B0(n117), .Y(n119) );
  OAI221X1 U6 ( .A0(addr[2]), .A1(n80), .B0(n118), .B1(n105), .C0(n79), .Y(
        dout[1]) );
  INVX4 U7 ( .A(addr[5]), .Y(n12) );
  OAI31X1 U8 ( .A0(n108), .A1(addr[5]), .A2(n6), .B0(n107), .Y(n109) );
  AOI222XL U9 ( .A0(n16), .A1(n72), .B0(n113), .B1(n7), .C0(addr[1]), .C1(n71), 
        .Y(n114) );
  OAI222X1 U10 ( .A0(addr[1]), .A1(n84), .B0(n85), .B1(n74), .C0(n71), .C1(
        n107), .Y(n75) );
  NAND2XL U11 ( .A(n1), .B(addr[5]), .Y(n84) );
  AOI211XL U13 ( .A0(n83), .A1(n12), .B0(n82), .C0(n8), .Y(n92) );
  NAND2XL U14 ( .A(n16), .B(n12), .Y(n74) );
  CLKINVX1 U15 ( .A(n118), .Y(n5) );
  CLKINVX1 U16 ( .A(n115), .Y(n15) );
  CLKINVX1 U17 ( .A(n112), .Y(n3) );
  OAI21X1 U18 ( .A0(n10), .A1(n6), .B0(n4), .Y(n112) );
  AOI22X1 U19 ( .A0(n11), .A1(n111), .B0(n6), .B1(n113), .Y(n93) );
  OAI211X1 U21 ( .A0(n7), .A1(n115), .B0(n93), .C0(n9), .Y(n94) );
  CLKINVX1 U22 ( .A(n85), .Y(n11) );
  NAND2X1 U23 ( .A(n97), .B(n71), .Y(n105) );
  NAND2X1 U24 ( .A(n113), .B(n5), .Y(n98) );
  NAND2X1 U25 ( .A(n10), .B(n97), .Y(n107) );
  NAND2X1 U26 ( .A(n118), .B(n85), .Y(n110) );
  OAI21XL U27 ( .A0(n15), .A1(n12), .B0(n108), .Y(n95) );
  CLKINVX1 U28 ( .A(n84), .Y(n14) );
  CLKINVX1 U29 ( .A(addr[2]), .Y(n4) );
  OAI31X1 U30 ( .A0(n16), .A1(addr[6]), .A2(n12), .B0(n87), .Y(n88) );
  OAI21XL U31 ( .A0(n113), .A1(n13), .B0(n11), .Y(n87) );
  OAI211X1 U32 ( .A0(n76), .A1(n16), .B0(n98), .C0(n9), .Y(n77) );
  AOI222XL U35 ( .A0(addr[5]), .A1(addr[6]), .B0(n111), .B1(addr[1]), .C0(n6), 
        .C1(n2), .Y(n76) );
  NAND3XL U36 ( .A(n11), .B(n71), .C(addr[4]), .Y(n117) );
  OAI22XL U37 ( .A0(n116), .A1(n115), .B0(n1), .B1(n112), .Y(n78) );
  CLKINVX3 U38 ( .A(addr[4]), .Y(n16) );
  OAI2BB2XL U39 ( .B0(n115), .B1(n106), .A0N(n12), .A1N(n86), .Y(n89) );
  OAI221XL U40 ( .A0(n116), .A1(addr[4]), .B0(n108), .B1(addr[1]), .C0(n117), 
        .Y(n86) );
  CLKINVX1 U41 ( .A(addr[6]), .Y(n72) );
  CLKINVX1 U42 ( .A(n81), .Y(n8) );
  OAI21XL U44 ( .A0(n96), .A1(n118), .B0(n93), .Y(n82) );
  NAND3X1 U46 ( .A(n101), .B(n100), .C(n99), .Y(n102) );
  AOI32X1 U47 ( .A0(n96), .A1(n71), .A2(n10), .B0(n11), .B1(n95), .Y(n101) );
  AOI2BB2XL U48 ( .B0(n7), .B1(n121), .A0N(n98), .A1N(addr[5]), .Y(n99) );
  OAI21XL U49 ( .A0(n97), .A1(n13), .B0(n6), .Y(n100) );
  AOI2BB2XL U50 ( .B0(n6), .B1(n123), .A0N(n122), .A1N(n4), .Y(n124) );
  AOI211XL U59 ( .A0(n6), .A1(n121), .B0(n120), .C0(n119), .Y(n122) );
  OAI22XL U60 ( .A0(n116), .A1(n115), .B0(addr[5]), .B1(n114), .Y(n120) );
  CLKINVX1 U61 ( .A(n75), .Y(n9) );
  AOI32XL U62 ( .A0(n10), .A1(n96), .A2(n1), .B0(addr[1]), .B1(n121), .Y(n81)
         );
  OAI211X1 U63 ( .A0(addr[2]), .A1(n126), .B0(n125), .C0(n124), .Y(dout[4]) );
  AOI32X1 U64 ( .A0(n11), .A1(n13), .A2(n2), .B0(n3), .B1(n14), .Y(n125) );
  AOI221XL U65 ( .A0(n5), .A1(n111), .B0(n15), .B1(n110), .C0(n109), .Y(n126)
         );
  AOI222XL U66 ( .A0(n6), .A1(n13), .B0(n121), .B1(n116), .C0(n2), .C1(n73), 
        .Y(n80) );
  AOI22XL U67 ( .A0(n78), .A1(n12), .B0(addr[2]), .B1(n77), .Y(n79) );
  OAI211X1 U68 ( .A0(n106), .A1(n105), .B0(n104), .C0(n103), .Y(dout[3]) );
  AOI32X1 U69 ( .A0(n2), .A1(n13), .A2(n10), .B0(n94), .B1(n4), .Y(n104) );
  AOI22XL U70 ( .A0(addr[2]), .A1(n102), .B0(n5), .B1(n123), .Y(n103) );
  NAND2XL U71 ( .A(n111), .B(addr[4]), .Y(n91) );
  AOI211X1 U72 ( .A0(n14), .A1(n110), .B0(n89), .C0(n88), .Y(n90) );
  CLKINVX3 U73 ( .A(n106), .Y(n6) );
  CLKINVX3 U74 ( .A(addr[1]), .Y(n7) );
  CLKINVX3 U75 ( .A(n96), .Y(n13) );
  CLKINVX3 U76 ( .A(n2), .Y(n71) );
endmodule


module sbox5_1 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121;

  OAI222X4 U18 ( .A0(addr[3]), .A1(n106), .B0(n8), .B1(n90), .C0(n13), .C1(n16), .Y(n93) );
  OAI22X2 U40 ( .A0(addr[5]), .A1(n106), .B0(n68), .B1(n114), .Y(n116) );
  NOR2X2 U41 ( .A(n3), .B(addr[3]), .Y(n102) );
  NAND2X2 U45 ( .A(addr[6]), .B(n16), .Y(n114) );
  NAND2X2 U50 ( .A(n16), .B(n8), .Y(n110) );
  NAND2X2 U52 ( .A(addr[1]), .B(n8), .Y(n113) );
  NAND2X2 U54 ( .A(addr[1]), .B(addr[6]), .Y(n106) );
  NAND2X2 U55 ( .A(addr[3]), .B(n13), .Y(n121) );
  OAI221X4 U1 ( .A0(n111), .A1(n110), .B0(n121), .B1(n114), .C0(n109), .Y(n112) );
  OAI221X4 U2 ( .A0(n107), .A1(n121), .B0(n111), .B1(n113), .C0(n85), .Y(n86)
         );
  OAI31X1 U3 ( .A0(n69), .A1(addr[5]), .A2(addr[1]), .B0(n81), .Y(n73) );
  CLKINVX1 U4 ( .A(addr[5]), .Y(n1) );
  OAI221X4 U5 ( .A0(n13), .A1(n114), .B0(n68), .B1(n113), .C0(n120), .Y(n115)
         );
  AOI221XL U6 ( .A0(n93), .A1(n1), .B0(n9), .B1(n14), .C0(n92), .Y(n105) );
  INVX3 U7 ( .A(addr[5]), .Y(n68) );
  OAI32X1 U8 ( .A0(n114), .A1(addr[5]), .A2(n3), .B0(n12), .B1(n107), .Y(n79)
         );
  AOI32XL U9 ( .A0(n14), .A1(n98), .A2(n7), .B0(n2), .B1(n73), .Y(n77) );
  CLKBUFX3 U10 ( .A(addr[4]), .Y(n2) );
  CLKINVX1 U11 ( .A(n81), .Y(n10) );
  NAND2X1 U12 ( .A(n11), .B(n14), .Y(n81) );
  CLKINVX1 U13 ( .A(n110), .Y(n5) );
  CLKXOR2X2 U14 ( .A(n69), .B(n68), .Y(n94) );
  AOI2BB1X1 U15 ( .A0N(n13), .A1N(n1), .B0(n14), .Y(n111) );
  NOR2X1 U16 ( .A(n121), .B(n68), .Y(n91) );
  NOR2BX1 U17 ( .AN(n116), .B(n90), .Y(n83) );
  NAND2X1 U19 ( .A(n5), .B(n68), .Y(n120) );
  CLKINVX1 U20 ( .A(n113), .Y(n7) );
  NAND2X1 U21 ( .A(n7), .B(n68), .Y(n107) );
  CLKINVX1 U22 ( .A(n121), .Y(n12) );
  OAI31X1 U23 ( .A0(n70), .A1(n14), .A2(n113), .B0(n99), .Y(n72) );
  CLKINVX1 U24 ( .A(n106), .Y(n9) );
  OAI2BB2XL U25 ( .B0(n1), .B1(n113), .A0N(n98), .A1N(n11), .Y(n101) );
  CLKINVX1 U26 ( .A(n114), .Y(n11) );
  CLKINVX1 U27 ( .A(n90), .Y(n15) );
  CLKINVX1 U28 ( .A(addr[1]), .Y(n16) );
  CLKINVX1 U29 ( .A(addr[3]), .Y(n69) );
  CLKINVX1 U30 ( .A(addr[6]), .Y(n8) );
  AOI211X1 U31 ( .A0(n91), .A1(addr[1]), .B0(n80), .C0(n79), .Y(n89) );
  OAI2BB2XL U32 ( .B0(n111), .B1(n106), .A0N(n94), .A1N(n5), .Y(n80) );
  AOI211X1 U33 ( .A0(n102), .A1(n84), .B0(n83), .C0(n82), .Y(n85) );
  OAI21XL U34 ( .A0(n8), .A1(n1), .B0(n106), .Y(n84) );
  NOR3XL U35 ( .A(n94), .B(n3), .C(n110), .Y(n82) );
  AOI222XL U36 ( .A0(n9), .A1(n15), .B0(addr[5]), .B1(n108), .C0(n6), .C1(n13), 
        .Y(n109) );
  CLKINVX1 U37 ( .A(n107), .Y(n6) );
  OAI21XL U38 ( .A0(addr[6]), .A1(addr[3]), .B0(n106), .Y(n108) );
  NAND2X1 U39 ( .A(addr[3]), .B(n3), .Y(n90) );
  NAND2X1 U42 ( .A(n2), .B(addr[5]), .Y(n98) );
  NAND2X1 U43 ( .A(n3), .B(n69), .Y(n97) );
  OAI21XL U44 ( .A0(addr[1]), .A1(n97), .B0(n96), .Y(n103) );
  AOI33XL U46 ( .A0(n3), .A1(n95), .A2(addr[5]), .B0(n94), .B1(n13), .B2(
        addr[1]), .Y(n96) );
  OAI21XL U47 ( .A0(n16), .A1(n69), .B0(n114), .Y(n95) );
  OAI21XL U48 ( .A0(addr[6]), .A1(n121), .B0(n99), .Y(n100) );
  NAND2X1 U49 ( .A(n71), .B(n5), .Y(n99) );
  XOR2X1 U51 ( .A(n70), .B(n3), .Y(n71) );
  AOI2BB2XL U53 ( .B0(n102), .B1(n116), .A0N(n2), .A1N(n75), .Y(n76) );
  AOI211X1 U56 ( .A0(n4), .A1(n3), .B0(n74), .C0(n83), .Y(n75) );
  AO22XL U57 ( .A0(n7), .A1(n12), .B0(addr[6]), .B1(n102), .Y(n74) );
  CLKINVX1 U58 ( .A(n120), .Y(n4) );
  CLKINVX1 U59 ( .A(n2), .Y(n70) );
  AO22XL U60 ( .A0(n7), .A1(n15), .B0(addr[6]), .B1(n91), .Y(n92) );
  AOI222XL U61 ( .A0(n116), .A1(n13), .B0(addr[3]), .B1(n115), .C0(n7), .C1(
        n14), .Y(n117) );
  OAI221X1 U62 ( .A0(n2), .A1(n105), .B0(n110), .B1(n121), .C0(n104), .Y(
        dout[3]) );
  AOI222XL U63 ( .A0(n2), .A1(n103), .B0(n102), .B1(n101), .C0(n100), .C1(n1), 
        .Y(n104) );
  OAI211X1 U64 ( .A0(n121), .A1(n120), .B0(n119), .C0(n118), .Y(dout[4]) );
  AOI32XL U65 ( .A0(n14), .A1(n114), .A2(addr[5]), .B0(n2), .B1(n112), .Y(n119) );
  AOI2BB2X1 U66 ( .B0(n10), .B1(n68), .A0N(n2), .A1N(n117), .Y(n118) );
  OAI211X1 U67 ( .A0(n2), .A1(n89), .B0(n88), .C0(n87), .Y(dout[2]) );
  AOI33XL U68 ( .A0(n12), .A1(n98), .A2(n11), .B0(n3), .B1(n94), .B2(n5), .Y(
        n88) );
  AOI222XL U69 ( .A0(n10), .A1(n68), .B0(n2), .B1(n86), .C0(n91), .C1(n9), .Y(
        n87) );
  OAI211X1 U70 ( .A0(n78), .A1(n68), .B0(n77), .C0(n76), .Y(dout[1]) );
  AOI221XL U71 ( .A0(n12), .A1(addr[1]), .B0(n9), .B1(n14), .C0(n72), .Y(n78)
         );
  BUFX4 U72 ( .A(addr[2]), .Y(n3) );
  CLKINVX3 U73 ( .A(n3), .Y(n13) );
  CLKINVX3 U74 ( .A(n97), .Y(n14) );
endmodule


module sbox6_1 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147;

  NAND2X2 U39 ( .A(n138), .B(addr[3]), .Y(n147) );
  NOR2X2 U47 ( .A(n83), .B(n81), .Y(n138) );
  NOR2X2 U50 ( .A(n10), .B(n4), .Y(n119) );
  NOR2X2 U58 ( .A(n85), .B(n10), .Y(n125) );
  NAND2X2 U61 ( .A(n97), .B(n103), .Y(n112) );
  NOR2X2 U62 ( .A(n17), .B(addr[1]), .Y(n103) );
  NOR2X2 U63 ( .A(n85), .B(addr[3]), .Y(n97) );
  NAND2X2 U64 ( .A(n117), .B(n131), .Y(n140) );
  NOR2X2 U65 ( .A(n5), .B(addr[3]), .Y(n131) );
  NOR2X2 U66 ( .A(n84), .B(addr[6]), .Y(n117) );
  NOR2X1 U1 ( .A(n83), .B(addr[3]), .Y(n102) );
  OAI222X1 U2 ( .A0(n91), .A1(n12), .B0(n3), .B1(n11), .C0(addr[5]), .C1(n8), 
        .Y(n92) );
  CLKINVX1 U3 ( .A(addr[3]), .Y(n1) );
  INVX3 U4 ( .A(addr[3]), .Y(n10) );
  CLKINVX1 U5 ( .A(n85), .Y(n2) );
  INVX4 U6 ( .A(n4), .Y(n85) );
  CLKBUFX3 U7 ( .A(addr[4]), .Y(n4) );
  CLKINVX1 U8 ( .A(n83), .Y(n3) );
  BUFX4 U9 ( .A(addr[2]), .Y(n5) );
  OAI221X1 U10 ( .A0(n17), .A1(n9), .B0(n10), .B1(n14), .C0(n86), .Y(n90) );
  INVX2 U11 ( .A(n96), .Y(n14) );
  NOR2X4 U12 ( .A(addr[1]), .B(addr[6]), .Y(n130) );
  OAI22X1 U13 ( .A0(n10), .A1(n17), .B0(addr[1]), .B1(n8), .Y(n142) );
  OAI221X4 U14 ( .A0(n123), .A1(n16), .B0(n81), .B1(n12), .C0(n13), .Y(n124)
         );
  NOR2X4 U15 ( .A(n5), .B(addr[5]), .Y(n143) );
  INVX1 U16 ( .A(n130), .Y(n82) );
  CLKINVX1 U17 ( .A(n125), .Y(n9) );
  NAND2X1 U18 ( .A(n82), .B(n14), .Y(n105) );
  INVXL U19 ( .A(n121), .Y(n6) );
  CLKINVX1 U20 ( .A(n138), .Y(n18) );
  AOI211X1 U21 ( .A0(n12), .A1(n10), .B0(n131), .C0(n143), .Y(n121) );
  CLKINVX1 U22 ( .A(n117), .Y(n81) );
  CLKINVX1 U23 ( .A(n119), .Y(n8) );
  NOR2X1 U24 ( .A(n14), .B(n123), .Y(n144) );
  NOR2X1 U25 ( .A(n84), .B(n17), .Y(n96) );
  CLKINVX1 U26 ( .A(n103), .Y(n16) );
  OAI211X1 U27 ( .A0(n82), .A1(n9), .B0(n104), .C0(n112), .Y(n108) );
  OAI21XL U28 ( .A0(n103), .A1(n117), .B0(n102), .Y(n104) );
  OAI21XL U29 ( .A0(n132), .A1(n17), .B0(n1), .Y(n86) );
  AOI21X1 U30 ( .A0(n85), .A1(n102), .B0(n125), .Y(n91) );
  OAI2BB2XL U31 ( .B0(n143), .B1(n82), .A0N(n143), .A1N(n117), .Y(n118) );
  CLKINVX1 U32 ( .A(n122), .Y(n13) );
  CLKINVX1 U33 ( .A(n126), .Y(n15) );
  CLKINVX1 U34 ( .A(n97), .Y(n11) );
  NAND2BX1 U35 ( .AN(n144), .B(n137), .Y(n107) );
  CLKINVX1 U36 ( .A(addr[1]), .Y(n84) );
  NOR2X1 U37 ( .A(n14), .B(n3), .Y(n122) );
  NOR2X1 U38 ( .A(addr[1]), .B(n2), .Y(n132) );
  OAI22X1 U40 ( .A0(n8), .A1(n81), .B0(n5), .B1(n15), .Y(n88) );
  NAND2X1 U41 ( .A(n5), .B(n12), .Y(n123) );
  NAND4X1 U42 ( .A(n147), .B(n140), .C(n100), .D(n99), .Y(n101) );
  AOI222XL U43 ( .A0(n98), .A1(n83), .B0(n102), .B1(n130), .C0(n97), .C1(n105), 
        .Y(n99) );
  NAND3X1 U44 ( .A(n5), .B(n8), .C(n96), .Y(n100) );
  OAI221X1 U45 ( .A0(n10), .A1(n16), .B0(n8), .B1(n17), .C0(n15), .Y(n98) );
  AOI22X1 U46 ( .A0(n4), .A1(n115), .B0(addr[5]), .B1(n114), .Y(n129) );
  OAI21XL U48 ( .A0(n121), .A1(n82), .B0(n147), .Y(n115) );
  OAI21XL U49 ( .A0(n113), .A1(n83), .B0(n112), .Y(n114) );
  AOI221XL U51 ( .A0(n119), .A1(n84), .B0(n130), .B1(addr[3]), .C0(n111), .Y(
        n113) );
  OAI22XL U52 ( .A0(n81), .A1(n85), .B0(addr[3]), .B1(n14), .Y(n111) );
  AOI211X1 U53 ( .A0(n4), .A1(n135), .B0(n134), .C0(n133), .Y(n136) );
  OA21XL U54 ( .A0(n1), .A1(n3), .B0(n132), .Y(n133) );
  OAI2BB2XL U55 ( .B0(n2), .B1(n13), .A0N(n131), .A1N(n130), .Y(n134) );
  OAI22X1 U56 ( .A0(n5), .A1(n81), .B0(n83), .B1(n14), .Y(n135) );
  CLKINVX3 U57 ( .A(addr[5]), .Y(n12) );
  AOI2BB2X1 U59 ( .B0(n5), .B1(n130), .A0N(n3), .A1N(n16), .Y(n137) );
  NOR2X1 U60 ( .A(n16), .B(n2), .Y(n126) );
  AOI2BB2XL U67 ( .B0(n143), .B1(n90), .A0N(n89), .A1N(n12), .Y(n94) );
  AOI211X1 U68 ( .A0(n122), .A1(n4), .B0(n88), .C0(n87), .Y(n89) );
  OAI32X1 U69 ( .A0(n16), .A1(n10), .A2(n83), .B0(n18), .B1(n11), .Y(n87) );
  NAND3X1 U70 ( .A(n147), .B(n140), .C(n139), .Y(n141) );
  AOI32X1 U71 ( .A0(n5), .A1(n84), .A2(n4), .B0(n138), .B1(n85), .Y(n139) );
  AO22XL U72 ( .A0(n143), .A1(n2), .B0(n116), .B1(n85), .Y(n120) );
  OAI21XL U73 ( .A0(n3), .A1(n12), .B0(n123), .Y(n116) );
  CLKINVX1 U74 ( .A(n106), .Y(n7) );
  AOI32XL U75 ( .A0(n105), .A1(n85), .A2(n1), .B0(addr[1]), .B1(n125), .Y(n106) );
  OAI211X1 U76 ( .A0(n2), .A1(n147), .B0(n146), .C0(n145), .Y(dout[4]) );
  AOI222XL U77 ( .A0(n144), .A1(n10), .B0(n143), .B1(n142), .C0(n141), .C1(n12), .Y(n145) );
  OA22X1 U78 ( .A0(n9), .A1(n137), .B0(n136), .B1(n12), .Y(n146) );
  NAND3X1 U79 ( .A(n129), .B(n128), .C(n127), .Y(dout[3]) );
  AOI32XL U80 ( .A0(n120), .A1(n10), .A2(addr[1]), .B0(n119), .B1(n118), .Y(
        n128) );
  AOI222XL U81 ( .A0(n144), .A1(n85), .B0(n126), .B1(n6), .C0(n125), .C1(n124), 
        .Y(n127) );
  NAND3BX1 U82 ( .AN(n95), .B(n94), .C(n93), .Y(dout[1]) );
  OAI222X1 U83 ( .A0(n140), .A1(n4), .B0(n112), .B1(n83), .C0(n14), .C1(n91), 
        .Y(n95) );
  AOI32XL U84 ( .A0(addr[1]), .A1(n12), .A2(n125), .B0(n130), .B1(n92), .Y(n93) );
  OAI211X1 U85 ( .A0(n85), .A1(n140), .B0(n110), .C0(n109), .Y(dout[2]) );
  AOI222XL U86 ( .A0(n108), .A1(n12), .B0(n143), .B1(n7), .C0(n119), .C1(n107), 
        .Y(n109) );
  AOI2BB2XL U87 ( .B0(addr[5]), .B1(n101), .A0N(n83), .A1N(n112), .Y(n110) );
  CLKINVX3 U88 ( .A(addr[6]), .Y(n17) );
  CLKINVX3 U89 ( .A(n5), .Y(n83) );
endmodule


module sbox7_1 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148;

  OAI222X4 U19 ( .A0(n19), .A1(n129), .B0(n4), .B1(n15), .C0(addr[1]), .C1(n7), 
        .Y(n122) );
  OAI33X4 U33 ( .A0(addr[1]), .A1(n4), .A2(n5), .B0(n16), .B1(n86), .B2(n13), 
        .Y(n97) );
  NOR2X2 U44 ( .A(n87), .B(n4), .Y(n116) );
  NOR2X2 U48 ( .A(addr[1]), .B(addr[6]), .Y(n136) );
  NOR2X2 U51 ( .A(n83), .B(n87), .Y(n125) );
  NOR2X2 U52 ( .A(n16), .B(addr[3]), .Y(n131) );
  NOR2X2 U58 ( .A(n93), .B(n124), .Y(n142) );
  NOR2X2 U60 ( .A(n85), .B(addr[1]), .Y(n93) );
  NOR2X2 U62 ( .A(n11), .B(n3), .Y(n137) );
  NOR2X2 U65 ( .A(n85), .B(n17), .Y(n140) );
  NAND2X1 U1 ( .A(n3), .B(n4), .Y(n119) );
  CLKBUFX3 U2 ( .A(addr[4]), .Y(n4) );
  CLKINVX1 U3 ( .A(n11), .Y(n1) );
  CLKINVX1 U4 ( .A(n86), .Y(n2) );
  CLKBUFX3 U5 ( .A(addr[2]), .Y(n5) );
  OAI31X1 U6 ( .A0(n87), .A1(n11), .A2(n17), .B0(n117), .Y(n121) );
  NOR2X4 U7 ( .A(n17), .B(addr[6]), .Y(n124) );
  OAI22X1 U8 ( .A0(addr[1]), .A1(n7), .B0(n5), .B1(n113), .Y(n100) );
  OAI22X1 U9 ( .A0(n4), .A1(n83), .B0(addr[3]), .B1(n10), .Y(n103) );
  AOI211XL U10 ( .A0(n2), .A1(n14), .B0(n131), .C0(n130), .Y(n132) );
  NOR3XL U11 ( .A(n19), .B(addr[3]), .C(n2), .Y(n130) );
  OAI21XL U12 ( .A0(n3), .A1(n1), .B0(n119), .Y(n89) );
  BUFX4 U13 ( .A(addr[5]), .Y(n3) );
  AOI221XL U14 ( .A0(n140), .A1(n89), .B0(n109), .B1(n14), .C0(n88), .Y(n96)
         );
  CLKINVX1 U15 ( .A(n140), .Y(n16) );
  OAI2BB2XL U16 ( .B0(n142), .B1(n10), .A0N(n141), .A1N(n140), .Y(n143) );
  CLKINVX1 U17 ( .A(n125), .Y(n21) );
  CLKINVX1 U18 ( .A(n142), .Y(n14) );
  NAND2X1 U20 ( .A(n21), .B(n84), .Y(n105) );
  CLKINVX1 U21 ( .A(n123), .Y(n6) );
  CLKINVX1 U22 ( .A(n109), .Y(n9) );
  NAND2X1 U23 ( .A(n124), .B(n87), .Y(n113) );
  CLKINVX1 U24 ( .A(n137), .Y(n10) );
  NOR2X1 U25 ( .A(n10), .B(n87), .Y(n109) );
  CLKINVX1 U26 ( .A(n136), .Y(n19) );
  OAI22XL U27 ( .A0(n137), .A1(n15), .B0(n17), .B1(n9), .Y(n146) );
  OAI21X1 U28 ( .A0(n11), .A1(n21), .B0(n129), .Y(n141) );
  NAND2X1 U29 ( .A(n116), .B(n83), .Y(n129) );
  CLKINVX1 U30 ( .A(n93), .Y(n18) );
  OAI21XL U31 ( .A0(n119), .A1(n18), .B0(n118), .Y(n120) );
  OAI21XL U32 ( .A0(n125), .A1(n137), .B0(n124), .Y(n118) );
  NOR2X1 U34 ( .A(n83), .B(n7), .Y(n123) );
  CLKINVX1 U35 ( .A(n145), .Y(n7) );
  OAI22XL U36 ( .A0(n137), .A1(n113), .B0(n85), .B1(n6), .Y(n88) );
  CLKINVX1 U37 ( .A(n116), .Y(n13) );
  CLKINVX1 U38 ( .A(n131), .Y(n15) );
  CLKINVX1 U39 ( .A(n134), .Y(n84) );
  NOR2XL U40 ( .A(n125), .B(n11), .Y(n110) );
  CLKINVX1 U41 ( .A(n119), .Y(n12) );
  CLKINVX1 U42 ( .A(n103), .Y(n8) );
  OA21XL U43 ( .A0(n20), .A1(n18), .B0(n117), .Y(n102) );
  CLKINVX1 U45 ( .A(n105), .Y(n20) );
  OAI2BB1XL U46 ( .A0N(n103), .A1N(n124), .B0(n102), .Y(n104) );
  OAI22X1 U47 ( .A0(n83), .A1(n13), .B0(n4), .B1(n84), .Y(n112) );
  NOR4X1 U49 ( .A(n4), .B(addr[3]), .C(n17), .D(n86), .Y(n99) );
  XNOR2X1 U50 ( .A(addr[6]), .B(n5), .Y(n101) );
  AOI211X1 U53 ( .A0(n116), .A1(addr[6]), .B0(n115), .C0(n114), .Y(n128) );
  OAI222X1 U54 ( .A0(n111), .A1(n16), .B0(n110), .B1(n18), .C0(n19), .C1(n9), 
        .Y(n115) );
  OAI2BB2XL U55 ( .B0(n12), .B1(n113), .A0N(n17), .A1N(n112), .Y(n114) );
  OA21XL U56 ( .A0(n87), .A1(n3), .B0(n6), .Y(n111) );
  NAND2X1 U57 ( .A(n5), .B(n136), .Y(n133) );
  CLKINVX1 U59 ( .A(addr[6]), .Y(n85) );
  AOI211X1 U61 ( .A0(n131), .A1(n3), .B0(n92), .C0(n91), .Y(n95) );
  OAI221X1 U63 ( .A0(n17), .A1(n7), .B0(n16), .B1(n10), .C0(n102), .Y(n92) );
  OAI31X1 U64 ( .A0(n87), .A1(n11), .A2(n19), .B0(n90), .Y(n91) );
  AO21XL U66 ( .A0(n119), .A1(n129), .B0(addr[6]), .Y(n90) );
  NOR2X1 U67 ( .A(n11), .B(addr[3]), .Y(n145) );
  AOI21XL U68 ( .A0(addr[3]), .A1(n98), .B0(n97), .Y(n108) );
  OAI2BB1XL U69 ( .A0N(n86), .A1N(n124), .B0(n133), .Y(n98) );
  NAND3X1 U70 ( .A(n136), .B(n87), .C(n3), .Y(n117) );
  NOR2X1 U71 ( .A(addr[3]), .B(n3), .Y(n134) );
  OAI21X1 U72 ( .A0(n5), .A1(n142), .B0(n133), .Y(n138) );
  OAI22XL U73 ( .A0(n142), .A1(n13), .B0(n1), .B1(n132), .Y(n135) );
  AO21X1 U74 ( .A0(n139), .A1(n83), .B0(n138), .Y(n144) );
  OAI21XL U75 ( .A0(n2), .A1(n17), .B0(n18), .Y(n139) );
  OAI221X1 U76 ( .A0(n3), .A1(n108), .B0(n107), .B1(n83), .C0(n106), .Y(
        dout[2]) );
  AOI32X1 U77 ( .A0(n105), .A1(n86), .A2(n140), .B0(n5), .B1(n104), .Y(n106)
         );
  AOI211X1 U78 ( .A0(n101), .A1(n4), .B0(n100), .C0(n99), .Y(n107) );
  OAI211X1 U79 ( .A0(n128), .A1(n86), .B0(n127), .C0(n126), .Y(dout[3]) );
  AOI32XL U80 ( .A0(n125), .A1(n1), .A2(n124), .B0(n123), .B1(n136), .Y(n126)
         );
  OAI31X1 U81 ( .A0(n122), .A1(n121), .A2(n120), .B0(n86), .Y(n127) );
  NAND2X1 U82 ( .A(n148), .B(n147), .Y(dout[4]) );
  AOI222XL U83 ( .A0(n136), .A1(n141), .B0(n3), .B1(n135), .C0(n134), .C1(n138), .Y(n148) );
  AOI222XL U84 ( .A0(n5), .A1(n146), .B0(n145), .B1(n144), .C0(n143), .C1(n86), 
        .Y(n147) );
  OAI221X1 U85 ( .A0(n96), .A1(n86), .B0(n5), .B1(n95), .C0(n94), .Y(dout[1])
         );
  AOI2BB2X1 U86 ( .B0(n93), .B1(n112), .A0N(n133), .A1N(n8), .Y(n94) );
  CLKINVX3 U87 ( .A(n4), .Y(n11) );
  CLKINVX3 U88 ( .A(addr[1]), .Y(n17) );
  CLKINVX3 U89 ( .A(n3), .Y(n83) );
  CLKINVX3 U90 ( .A(n5), .Y(n86) );
  CLKINVX3 U91 ( .A(addr[3]), .Y(n87) );
endmodule


module sbox8_1 ( addr, dout );
  input [1:6] addr;
  output [1:4] dout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132;

  NAND2X2 U41 ( .A(addr[6]), .B(n74), .Y(n131) );
  NAND2X2 U48 ( .A(addr[4]), .B(n7), .Y(n123) );
  NAND2X2 U49 ( .A(n2), .B(n4), .Y(n87) );
  NAND2X2 U50 ( .A(addr[1]), .B(n14), .Y(n124) );
  NAND2X2 U54 ( .A(addr[2]), .B(n75), .Y(n116) );
  NAND2X2 U60 ( .A(addr[6]), .B(addr[1]), .Y(n105) );
  NAND2X2 U61 ( .A(n74), .B(n14), .Y(n108) );
  OAI32X1 U1 ( .A0(n14), .A1(addr[4]), .A2(n92), .B0(n115), .B1(n108), .Y(n96)
         );
  OAI31X1 U2 ( .A0(n123), .A1(addr[6]), .A2(n116), .B0(n109), .Y(n110) );
  OAI221X1 U3 ( .A0(n105), .A1(n87), .B0(addr[4]), .B1(n108), .C0(n86), .Y(n90) );
  NAND2X4 U4 ( .A(addr[4]), .B(n2), .Y(n115) );
  AOI222X1 U5 ( .A0(n88), .A1(addr[2]), .B0(n4), .B1(n8), .C0(n9), .C1(n92), 
        .Y(n114) );
  OAI222X1 U6 ( .A0(addr[2]), .A1(n126), .B0(n7), .B1(n125), .C0(n124), .C1(
        n123), .Y(n127) );
  AOI32XL U7 ( .A0(n12), .A1(n10), .A2(n2), .B0(n13), .B1(n117), .Y(n130) );
  OA21XL U8 ( .A0(n9), .A1(n75), .B0(n121), .Y(n78) );
  INVXL U9 ( .A(n119), .Y(n5) );
  INVX3 U10 ( .A(n2), .Y(n7) );
  BUFX4 U11 ( .A(addr[3]), .Y(n2) );
  CLKBUFX3 U12 ( .A(addr[5]), .Y(n1) );
  CLKINVX1 U13 ( .A(n108), .Y(n13) );
  CLKINVX1 U14 ( .A(n107), .Y(n6) );
  CLKINVX1 U15 ( .A(n93), .Y(n3) );
  NAND2X1 U16 ( .A(n7), .B(n4), .Y(n93) );
  NAND2X1 U17 ( .A(n9), .B(n75), .Y(n121) );
  OAI21XL U18 ( .A0(n115), .A1(n75), .B0(n107), .Y(n77) );
  OAI21X1 U19 ( .A0(n4), .A1(n75), .B0(n123), .Y(n88) );
  OAI31XL U20 ( .A0(n115), .A1(n74), .A2(n116), .B0(n118), .Y(n94) );
  CLKINVX1 U21 ( .A(n131), .Y(n16) );
  NAND2X1 U22 ( .A(n10), .B(n7), .Y(n107) );
  OAI22XL U23 ( .A0(n116), .A1(n123), .B0(n10), .B1(n115), .Y(n117) );
  OAI22XL U24 ( .A0(n123), .A1(n108), .B0(n131), .B1(n93), .Y(n95) );
  OAI2BB2XL U25 ( .B0(n115), .B1(n131), .A0N(n88), .A1N(n15), .Y(n89) );
  AOI211XL U26 ( .A0(n108), .A1(n105), .B0(n4), .C0(n121), .Y(n85) );
  CLKINVX1 U27 ( .A(n124), .Y(n12) );
  OAI22XL U28 ( .A0(n10), .A1(n123), .B0(n78), .B1(n87), .Y(n81) );
  NAND2BX2 U29 ( .AN(n78), .B(n7), .Y(n120) );
  NAND2XL U30 ( .A(n115), .B(n93), .Y(n104) );
  OAI2BB2XL U31 ( .B0(n106), .B1(n105), .A0N(n104), .A1N(n12), .Y(n111) );
  NOR2BXL U32 ( .AN(n123), .B(n103), .Y(n106) );
  NAND3X1 U33 ( .A(n104), .B(n74), .C(n10), .Y(n84) );
  AO21X1 U34 ( .A0(n10), .A1(n15), .B0(n101), .Y(n102) );
  OAI33X1 U35 ( .A0(n14), .A1(n7), .A2(n100), .B0(n9), .B1(n103), .B2(n124), 
        .Y(n101) );
  OA22XL U36 ( .A0(n107), .A1(n131), .B0(n120), .B1(n124), .Y(n98) );
  CLKINVX1 U37 ( .A(n125), .Y(n11) );
  OAI21XL U38 ( .A0(n12), .A1(n16), .B0(addr[4]), .Y(n86) );
  NAND2X1 U39 ( .A(n1), .B(n9), .Y(n100) );
  OAI221X1 U40 ( .A0(n124), .A1(n121), .B0(addr[1]), .B1(n120), .C0(n5), .Y(
        n128) );
  OAI31XL U42 ( .A0(n9), .A1(n74), .A2(n7), .B0(n118), .Y(n119) );
  NAND2X1 U43 ( .A(n15), .B(addr[2]), .Y(n125) );
  NAND4XL U44 ( .A(n16), .B(n1), .C(n2), .D(addr[2]), .Y(n109) );
  NAND3X1 U45 ( .A(n10), .B(n14), .C(n2), .Y(n118) );
  OAI21XL U46 ( .A0(n1), .A1(n87), .B0(n114), .Y(n76) );
  OAI22XL U47 ( .A0(n108), .A1(n120), .B0(n79), .B1(n100), .Y(n80) );
  AOI221XL U51 ( .A0(n16), .A1(n7), .B0(n15), .B1(n2), .C0(n91), .Y(n79) );
  NOR2X1 U52 ( .A(n1), .B(n2), .Y(n103) );
  NOR2X1 U53 ( .A(n87), .B(addr[6]), .Y(n91) );
  NOR2X1 U55 ( .A(n7), .B(n1), .Y(n92) );
  CLKINVX1 U56 ( .A(n100), .Y(n8) );
  OA21XL U57 ( .A0(n1), .A1(n115), .B0(n120), .Y(n132) );
  AOI221XL U58 ( .A0(n13), .A1(n2), .B0(n15), .B1(addr[4]), .C0(n122), .Y(n126) );
  OAI22XL U59 ( .A0(n2), .A1(n74), .B0(addr[4]), .B1(n131), .Y(n122) );
  OAI211X1 U62 ( .A0(addr[2]), .A1(n99), .B0(n98), .C0(n97), .Y(dout[2]) );
  AOI221XL U63 ( .A0(addr[2]), .A1(n96), .B0(n1), .B1(n95), .C0(n94), .Y(n97)
         );
  AOI221XL U64 ( .A0(n91), .A1(n1), .B0(n90), .B1(n75), .C0(n89), .Y(n99) );
  OAI211X1 U65 ( .A0(n132), .A1(n131), .B0(n130), .C0(n129), .Y(dout[4]) );
  AOI222XL U66 ( .A0(n128), .A1(n4), .B0(n1), .B1(n127), .C0(n6), .C1(n15), 
        .Y(n129) );
  NAND4BX1 U67 ( .AN(n85), .B(n84), .C(n83), .D(n82), .Y(dout[1]) );
  AOI221XL U68 ( .A0(n16), .A1(n81), .B0(n3), .B1(n11), .C0(n80), .Y(n82) );
  AOI22X1 U69 ( .A0(n15), .A1(n77), .B0(n12), .B1(n76), .Y(n83) );
  OAI211X1 U70 ( .A0(addr[1]), .A1(n114), .B0(n113), .C0(n112), .Y(dout[3]) );
  AOI221XL U71 ( .A0(n111), .A1(n9), .B0(n6), .B1(n13), .C0(n110), .Y(n112) );
  AOI2BB2XL U72 ( .B0(n102), .B1(n4), .A0N(n115), .A1N(n125), .Y(n113) );
  CLKINVX3 U73 ( .A(addr[4]), .Y(n4) );
  CLKINVX3 U74 ( .A(addr[2]), .Y(n9) );
  CLKINVX3 U75 ( .A(n116), .Y(n10) );
  CLKINVX3 U76 ( .A(addr[6]), .Y(n14) );
  CLKINVX3 U77 ( .A(n105), .Y(n15) );
  CLKINVX3 U78 ( .A(addr[1]), .Y(n74) );
  CLKINVX3 U79 ( .A(n1), .Y(n75) );
endmodule


module crp_1 ( P, R, K_sub );
  output [1:32] P;
  input [1:32] R;
  input [1:48] K_sub;
  wire   n1;
  wire   [1:48] X;

  sbox1_1 u0 ( .addr(X[1:6]), .dout({P[9], P[17], P[23], P[31]}) );
  sbox2_1 u1 ( .addr({X[7], n1, X[9:12]}), .dout({P[13], P[28], P[2], P[18]})
         );
  sbox3_1 u2 ( .addr(X[13:18]), .dout({P[24], P[16], P[30], P[6]}) );
  sbox4_1 u3 ( .addr(X[19:24]), .dout({P[26], P[20], P[10], P[1]}) );
  sbox5_1 u4 ( .addr(X[25:30]), .dout({P[8], P[14], P[25], P[3]}) );
  sbox6_1 u5 ( .addr(X[31:36]), .dout({P[4], P[29], P[11], P[19]}) );
  sbox7_1 u6 ( .addr(X[37:42]), .dout({P[32], P[12], P[22], P[7]}) );
  sbox8_1 u7 ( .addr(X[43:48]), .dout({P[5], P[27], P[15], P[21]}) );
  XOR2X1 U1 ( .A(R[1]), .B(K_sub[2]), .Y(X[2]) );
  CLKXOR2X4 U2 ( .A(R[29]), .B(K_sub[42]), .Y(X[42]) );
  CLKXOR2X4 U3 ( .A(R[5]), .B(K_sub[6]), .Y(X[6]) );
  CLKXOR2X4 U4 ( .A(R[16]), .B(K_sub[25]), .Y(X[25]) );
  CLKXOR2X4 U5 ( .A(R[8]), .B(K_sub[11]), .Y(X[11]) );
  CLKXOR2X4 U6 ( .A(R[20]), .B(K_sub[31]), .Y(X[31]) );
  CLKXOR2X4 U7 ( .A(R[16]), .B(K_sub[23]), .Y(X[23]) );
  CLKXOR2X4 U8 ( .A(R[10]), .B(K_sub[15]), .Y(X[15]) );
  XNOR2X1 U9 ( .A(R[5]), .B(K_sub[8]), .Y(X[8]) );
  INVX3 U10 ( .A(X[8]), .Y(n1) );
  CLKXOR2X4 U11 ( .A(R[31]), .B(K_sub[46]), .Y(X[46]) );
  CLKXOR2X4 U12 ( .A(R[22]), .B(K_sub[33]), .Y(X[33]) );
  CLKXOR2X4 U13 ( .A(R[29]), .B(K_sub[44]), .Y(X[44]) );
  CLKXOR2X4 U14 ( .A(R[12]), .B(K_sub[19]), .Y(X[19]) );
  CLKXOR2X4 U15 ( .A(R[26]), .B(K_sub[39]), .Y(X[39]) );
  CLKXOR2X4 U16 ( .A(R[20]), .B(K_sub[29]), .Y(X[29]) );
  CLKXOR2X2 U17 ( .A(R[4]), .B(K_sub[5]), .Y(X[5]) );
  CLKXOR2X2 U18 ( .A(R[15]), .B(K_sub[22]), .Y(X[22]) );
  CLKXOR2X2 U19 ( .A(R[24]), .B(K_sub[35]), .Y(X[35]) );
  CLKXOR2X2 U20 ( .A(R[21]), .B(K_sub[30]), .Y(X[30]) );
  CLKXOR2X2 U21 ( .A(R[12]), .B(K_sub[17]), .Y(X[17]) );
  CLKXOR2X2 U22 ( .A(R[32]), .B(K_sub[1]), .Y(X[1]) );
  CLKXOR2X2 U23 ( .A(R[13]), .B(K_sub[20]), .Y(X[20]) );
  CLKXOR2X2 U24 ( .A(R[18]), .B(K_sub[27]), .Y(X[27]) );
  CLKXOR2X2 U25 ( .A(R[8]), .B(K_sub[13]), .Y(X[13]) );
  CLKXOR2X2 U26 ( .A(R[4]), .B(K_sub[7]), .Y(X[7]) );
  CLKXOR2X2 U27 ( .A(R[24]), .B(K_sub[37]), .Y(X[37]) );
  CLKXOR2X2 U28 ( .A(R[28]), .B(K_sub[43]), .Y(X[43]) );
  CLKXOR2X2 U29 ( .A(R[1]), .B(K_sub[48]), .Y(X[48]) );
  CLKXOR2X2 U30 ( .A(R[17]), .B(K_sub[24]), .Y(X[24]) );
  CLKXOR2X2 U31 ( .A(R[9]), .B(K_sub[12]), .Y(X[12]) );
  CLKXOR2X2 U32 ( .A(R[13]), .B(K_sub[18]), .Y(X[18]) );
  CLKXOR2X2 U33 ( .A(R[25]), .B(K_sub[36]), .Y(X[36]) );
  XOR2X1 U34 ( .A(R[23]), .B(K_sub[34]), .Y(X[34]) );
  XOR2X1 U35 ( .A(R[9]), .B(K_sub[14]), .Y(X[14]) );
  XOR2X1 U36 ( .A(R[30]), .B(K_sub[45]), .Y(X[45]) );
  XOR2X1 U37 ( .A(R[21]), .B(K_sub[32]), .Y(X[32]) );
  XOR2X1 U38 ( .A(R[25]), .B(K_sub[38]), .Y(X[38]) );
  XOR2X1 U39 ( .A(R[27]), .B(K_sub[40]), .Y(X[40]) );
  XOR2X1 U40 ( .A(R[3]), .B(K_sub[4]), .Y(X[4]) );
  XOR2X1 U41 ( .A(R[11]), .B(K_sub[16]), .Y(X[16]) );
  XOR2X1 U42 ( .A(R[7]), .B(K_sub[10]), .Y(X[10]) );
  XOR2X1 U43 ( .A(R[14]), .B(K_sub[21]), .Y(X[21]) );
  XOR2X1 U44 ( .A(R[6]), .B(K_sub[9]), .Y(X[9]) );
  XOR2X1 U45 ( .A(R[2]), .B(K_sub[3]), .Y(X[3]) );
  XOR2X1 U46 ( .A(R[28]), .B(K_sub[41]), .Y(X[41]) );
  XOR2X1 U47 ( .A(R[17]), .B(K_sub[26]), .Y(X[26]) );
  XOR2X1 U48 ( .A(R[32]), .B(K_sub[47]), .Y(X[47]) );
  XOR2X1 U49 ( .A(R[19]), .B(K_sub[28]), .Y(X[28]) );
endmodule


module des ( desOut, desIn, key, decrypt, clk );
  output [63:0] desOut;
  input [63:0] desIn;
  input [55:0] key;
  input decrypt, clk;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85,
         N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99,
         N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132,
         N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176,
         N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187,
         N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198,
         N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N232, N233, N234, N235, N236, N237, N238, N239, N240, N241, N242,
         N243, N244, N245, N246, N247, N248, N249, N250, N251, N252, N253,
         N254, N255, N256, N257, N258, N259, N260, N261, N262, N263, N264,
         N265, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N364, N365, N366, N367, N368, N369, N370, N371, N372, N373, N374,
         N375, N376, N377, N378, N379, N380, N381, N382, N383, N384, N385,
         N386, N387, N388, N389, N390, N391, N392, N393, N394, N395, N396,
         N397, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N430, N431, N432, N433, N434, N435, N436, N437, N438, N439, N440,
         N441, N442, N443, N444, N445, N446, N447, N448, N449, N450, N451,
         N452, N453, N454, N455, N456, N457, N458, N459, N460, N461, N462,
         N463, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144;
  wire   [55:0] key_r;
  wire   [63:0] desIn_r;
  wire   [1:32] out15;
  wire   [1:32] L14;
  wire   [1:64] FP;
  wire   [1:48] K1;
  wire   [1:48] K2;
  wire   [1:48] K3;
  wire   [1:48] K4;
  wire   [1:48] K5;
  wire   [1:48] K6;
  wire   [1:48] K7;
  wire   [1:48] K8;
  wire   [1:48] K9;
  wire   [1:48] K10;
  wire   [1:48] K11;
  wire   [1:48] K12;
  wire   [1:48] K13;
  wire   [1:48] K14;
  wire   [1:48] K15;
  wire   [1:48] K16;
  wire   [1:32] out0;
  wire   [1:32] out1;
  wire   [1:32] R0;
  wire   [1:32] out2;
  wire   [1:32] R1;
  wire   [1:32] out3;
  wire   [1:32] R2;
  wire   [1:32] out4;
  wire   [1:32] R3;
  wire   [1:32] out5;
  wire   [1:32] R4;
  wire   [1:32] out6;
  wire   [1:32] R5;
  wire   [1:32] out7;
  wire   [1:32] R6;
  wire   [1:32] out8;
  wire   [1:32] R7;
  wire   [1:32] out9;
  wire   [1:32] R8;
  wire   [1:32] out10;
  wire   [1:32] R9;
  wire   [1:32] out11;
  wire   [1:32] R10;
  wire   [1:32] out12;
  wire   [1:32] R11;
  wire   [1:32] out13;
  wire   [1:32] R12;
  wire   [1:32] out14;
  wire   [1:32] R13;
  wire   [1:32] L0;
  wire   [1:32] L1;
  wire   [1:32] L2;
  wire   [1:32] L3;
  wire   [1:32] L4;
  wire   [1:32] L5;
  wire   [1:32] L6;
  wire   [1:32] L7;
  wire   [1:32] L8;
  wire   [1:32] L9;
  wire   [1:32] L10;
  wire   [1:32] L11;
  wire   [1:32] L12;
  wire   [1:32] L13;

  key_sel uk ( .clk(n120), .K(key_r), .decrypt(n1), .K1(K1), .K2(K2), .K3(K3), 
        .K4(K4), .K5(K5), .K6(K6), .K7(K7), .K8(K8), .K9(K9), .K10(K10), .K11(
        K11), .K12(K12), .K13(K13), .K14(K14), .K15(K15), .K16(K16) );
  crp_0 u0 ( .P(out0), .R({desIn_r[7], desIn_r[15], desIn_r[23], desIn_r[31], 
        desIn_r[39], desIn_r[47], desIn_r[55], desIn_r[63], desIn_r[5], 
        desIn_r[13], desIn_r[21], desIn_r[29], desIn_r[37], desIn_r[45], 
        desIn_r[53], desIn_r[61], desIn_r[3], desIn_r[11], desIn_r[19], 
        desIn_r[27], desIn_r[35], desIn_r[43], desIn_r[51], desIn_r[59], 
        desIn_r[1], desIn_r[9], desIn_r[17], desIn_r[25], desIn_r[33], 
        desIn_r[41], desIn_r[49], desIn_r[57]}), .K_sub(K1) );
  crp_15 u1 ( .P(out1), .R(R0), .K_sub(K2) );
  crp_14 u2 ( .P(out2), .R(R1), .K_sub(K3) );
  crp_13 u3 ( .P(out3), .R(R2), .K_sub(K4) );
  crp_12 u4 ( .P(out4), .R(R3), .K_sub(K5) );
  crp_11 u5 ( .P(out5), .R(R4), .K_sub(K6) );
  crp_10 u6 ( .P(out6), .R(R5), .K_sub(K7) );
  crp_9 u7 ( .P(out7), .R(R6), .K_sub(K8) );
  crp_8 u8 ( .P(out8), .R(R7), .K_sub(K9) );
  crp_7 u9 ( .P(out9), .R(R8), .K_sub(K10) );
  crp_6 u10 ( .P(out10), .R(R9), .K_sub(K11) );
  crp_5 u11 ( .P(out11), .R(R10), .K_sub(K12) );
  crp_4 u12 ( .P(out12), .R(R11), .K_sub(K13) );
  crp_3 u13 ( .P(out13), .R(R12), .K_sub(K14) );
  crp_2 u14 ( .P(out14), .R(R13), .K_sub(K15) );
  crp_1 u15 ( .P(out15), .R(FP[33:64]), .K_sub(K16) );
  DFFQX1 \desOut_reg[51]  ( .D(FP[55]), .CK(n138), .Q(desOut[51]) );
  DFFQX1 \desOut_reg[50]  ( .D(FP[23]), .CK(clk), .Q(desOut[50]) );
  DFFQX1 \desOut_reg[49]  ( .D(FP[63]), .CK(n137), .Q(desOut[49]) );
  DFFQX1 \desOut_reg[48]  ( .D(FP[31]), .CK(n136), .Q(desOut[48]) );
  DFFQX1 \desOut_reg[35]  ( .D(FP[53]), .CK(n109), .Q(desOut[35]) );
  DFFQX1 \desOut_reg[34]  ( .D(FP[21]), .CK(n110), .Q(desOut[34]) );
  DFFQX1 \desOut_reg[33]  ( .D(FP[61]), .CK(n111), .Q(desOut[33]) );
  DFFQX1 \desOut_reg[32]  ( .D(FP[29]), .CK(n86), .Q(desOut[32]) );
  DFFQX1 \desOut_reg[19]  ( .D(FP[51]), .CK(n123), .Q(desOut[19]) );
  DFFQX1 \desOut_reg[18]  ( .D(FP[19]), .CK(n124), .Q(desOut[18]) );
  DFFQX1 \desOut_reg[17]  ( .D(FP[59]), .CK(n125), .Q(desOut[17]) );
  DFFQX1 \desOut_reg[16]  ( .D(FP[27]), .CK(n126), .Q(desOut[16]) );
  DFFQX1 \desOut_reg[55]  ( .D(FP[39]), .CK(n139), .Q(desOut[55]) );
  DFFQX1 \desOut_reg[54]  ( .D(FP[7]), .CK(n136), .Q(desOut[54]) );
  DFFQX1 \desOut_reg[53]  ( .D(FP[47]), .CK(n135), .Q(desOut[53]) );
  DFFQX1 \desOut_reg[52]  ( .D(FP[15]), .CK(n134), .Q(desOut[52]) );
  DFFQX1 \desOut_reg[39]  ( .D(FP[37]), .CK(n112), .Q(desOut[39]) );
  DFFQX1 \desOut_reg[38]  ( .D(FP[5]), .CK(n113), .Q(desOut[38]) );
  DFFQX1 \desOut_reg[37]  ( .D(FP[45]), .CK(n114), .Q(desOut[37]) );
  DFFQX1 \desOut_reg[36]  ( .D(FP[13]), .CK(n115), .Q(desOut[36]) );
  DFFQX1 \desOut_reg[23]  ( .D(FP[35]), .CK(n87), .Q(desOut[23]) );
  DFFQX1 \desOut_reg[22]  ( .D(FP[3]), .CK(n127), .Q(desOut[22]) );
  DFFQX1 \desOut_reg[21]  ( .D(FP[43]), .CK(n8), .Q(desOut[21]) );
  DFFQX1 \desOut_reg[20]  ( .D(FP[11]), .CK(n53), .Q(desOut[20]) );
  DFFQX1 \desOut_reg[7]  ( .D(FP[33]), .CK(n122), .Q(desOut[7]) );
  DFFQX1 \desOut_reg[6]  ( .D(FP[1]), .CK(n112), .Q(desOut[6]) );
  DFFQX1 \desOut_reg[3]  ( .D(FP[49]), .CK(n121), .Q(desOut[3]) );
  DFFQX1 \desOut_reg[2]  ( .D(FP[17]), .CK(n122), .Q(desOut[2]) );
  DFFQX1 \desOut_reg[1]  ( .D(FP[57]), .CK(n111), .Q(desOut[1]) );
  DFFQX1 \desOut_reg[0]  ( .D(FP[25]), .CK(clk), .Q(desOut[0]) );
  DFFQX1 \desOut_reg[5]  ( .D(FP[41]), .CK(n47), .Q(desOut[5]) );
  DFFQX1 \desOut_reg[4]  ( .D(FP[9]), .CK(n117), .Q(desOut[4]) );
  DFFQX1 \desOut_reg[63]  ( .D(FP[40]), .CK(n131), .Q(desOut[63]) );
  DFFQX1 \desOut_reg[62]  ( .D(FP[8]), .CK(n130), .Q(desOut[62]) );
  DFFQX1 \desOut_reg[61]  ( .D(FP[48]), .CK(n141), .Q(desOut[61]) );
  DFFQX1 \desOut_reg[60]  ( .D(FP[16]), .CK(n117), .Q(desOut[60]) );
  DFFQX1 \desOut_reg[47]  ( .D(FP[38]), .CK(n129), .Q(desOut[47]) );
  DFFQX1 \desOut_reg[46]  ( .D(FP[6]), .CK(n128), .Q(desOut[46]) );
  DFFQX1 \desOut_reg[45]  ( .D(FP[46]), .CK(n81), .Q(desOut[45]) );
  DFFQX1 \desOut_reg[44]  ( .D(FP[14]), .CK(n28), .Q(desOut[44]) );
  DFFQX1 \desOut_reg[31]  ( .D(FP[36]), .CK(n103), .Q(desOut[31]) );
  DFFQX1 \desOut_reg[30]  ( .D(FP[4]), .CK(n128), .Q(desOut[30]) );
  DFFQX1 \desOut_reg[29]  ( .D(FP[44]), .CK(n80), .Q(desOut[29]) );
  DFFQX1 \desOut_reg[28]  ( .D(FP[12]), .CK(n105), .Q(desOut[28]) );
  DFFQX1 \desOut_reg[15]  ( .D(FP[34]), .CK(n143), .Q(desOut[15]) );
  DFFQX1 \desOut_reg[14]  ( .D(FP[2]), .CK(n135), .Q(desOut[14]) );
  DFFQX1 \desOut_reg[13]  ( .D(FP[42]), .CK(n95), .Q(desOut[13]) );
  DFFQX1 \desOut_reg[12]  ( .D(FP[10]), .CK(n98), .Q(desOut[12]) );
  DFFQX1 \desOut_reg[59]  ( .D(FP[56]), .CK(n133), .Q(desOut[59]) );
  DFFQX1 \desOut_reg[58]  ( .D(FP[24]), .CK(n140), .Q(desOut[58]) );
  DFFQX1 \desOut_reg[57]  ( .D(FP[64]), .CK(n132), .Q(desOut[57]) );
  DFFQX1 \desOut_reg[56]  ( .D(FP[32]), .CK(n98), .Q(desOut[56]) );
  DFFQX1 \desOut_reg[43]  ( .D(FP[54]), .CK(n118), .Q(desOut[43]) );
  DFFQX1 \desOut_reg[42]  ( .D(FP[22]), .CK(n138), .Q(desOut[42]) );
  DFFQX1 \desOut_reg[41]  ( .D(FP[62]), .CK(n116), .Q(desOut[41]) );
  DFFQX1 \desOut_reg[40]  ( .D(FP[30]), .CK(n103), .Q(desOut[40]) );
  DFFQX1 \desOut_reg[27]  ( .D(FP[52]), .CK(n106), .Q(desOut[27]) );
  DFFQX1 \desOut_reg[26]  ( .D(FP[20]), .CK(n107), .Q(desOut[26]) );
  DFFQX1 \desOut_reg[25]  ( .D(FP[60]), .CK(n108), .Q(desOut[25]) );
  DFFQX1 \desOut_reg[24]  ( .D(FP[28]), .CK(n104), .Q(desOut[24]) );
  DFFQX1 \desOut_reg[11]  ( .D(FP[50]), .CK(clk), .Q(desOut[11]) );
  DFFQX1 \desOut_reg[10]  ( .D(FP[18]), .CK(n137), .Q(desOut[10]) );
  DFFQX1 \desOut_reg[9]  ( .D(FP[58]), .CK(n144), .Q(desOut[9]) );
  DFFQX1 \desOut_reg[8]  ( .D(FP[26]), .CK(n144), .Q(desOut[8]) );
  DFFQX1 \desIn_r_reg[62]  ( .D(desIn[62]), .CK(n91), .Q(desIn_r[62]) );
  DFFQX1 \desIn_r_reg[60]  ( .D(desIn[60]), .CK(n90), .Q(desIn_r[60]) );
  DFFQX1 \desIn_r_reg[58]  ( .D(desIn[58]), .CK(n90), .Q(desIn_r[58]) );
  DFFQX1 \desIn_r_reg[56]  ( .D(desIn[56]), .CK(n90), .Q(desIn_r[56]) );
  DFFQX1 \desIn_r_reg[54]  ( .D(desIn[54]), .CK(n90), .Q(desIn_r[54]) );
  DFFQX1 \desIn_r_reg[52]  ( .D(desIn[52]), .CK(n89), .Q(desIn_r[52]) );
  DFFQX1 \desIn_r_reg[50]  ( .D(desIn[50]), .CK(n89), .Q(desIn_r[50]) );
  DFFQX1 \desIn_r_reg[48]  ( .D(desIn[48]), .CK(n89), .Q(desIn_r[48]) );
  DFFQX1 \desIn_r_reg[46]  ( .D(desIn[46]), .CK(n89), .Q(desIn_r[46]) );
  DFFQX1 \desIn_r_reg[44]  ( .D(desIn[44]), .CK(n89), .Q(desIn_r[44]) );
  DFFQX1 \desIn_r_reg[42]  ( .D(desIn[42]), .CK(n88), .Q(desIn_r[42]) );
  DFFQX1 \desIn_r_reg[40]  ( .D(desIn[40]), .CK(n88), .Q(desIn_r[40]) );
  DFFQX1 \desIn_r_reg[38]  ( .D(desIn[38]), .CK(n88), .Q(desIn_r[38]) );
  DFFQX1 \desIn_r_reg[36]  ( .D(desIn[36]), .CK(n88), .Q(desIn_r[36]) );
  DFFQX1 \desIn_r_reg[34]  ( .D(desIn[34]), .CK(n87), .Q(desIn_r[34]) );
  DFFQX1 \desIn_r_reg[32]  ( .D(desIn[32]), .CK(n87), .Q(desIn_r[32]) );
  DFFQX1 \desIn_r_reg[30]  ( .D(desIn[30]), .CK(n87), .Q(desIn_r[30]) );
  DFFQX1 \desIn_r_reg[28]  ( .D(desIn[28]), .CK(n87), .Q(desIn_r[28]) );
  DFFQX1 \desIn_r_reg[26]  ( .D(desIn[26]), .CK(n87), .Q(desIn_r[26]) );
  DFFQX1 \desIn_r_reg[24]  ( .D(desIn[24]), .CK(n86), .Q(desIn_r[24]) );
  DFFQX1 \desIn_r_reg[22]  ( .D(desIn[22]), .CK(n86), .Q(desIn_r[22]) );
  DFFQX1 \desIn_r_reg[20]  ( .D(desIn[20]), .CK(n86), .Q(desIn_r[20]) );
  DFFQX1 \desIn_r_reg[18]  ( .D(desIn[18]), .CK(n86), .Q(desIn_r[18]) );
  DFFQX1 \desIn_r_reg[16]  ( .D(desIn[16]), .CK(n85), .Q(desIn_r[16]) );
  DFFQX1 \desIn_r_reg[14]  ( .D(desIn[14]), .CK(n85), .Q(desIn_r[14]) );
  DFFQX1 \desIn_r_reg[12]  ( .D(desIn[12]), .CK(n85), .Q(desIn_r[12]) );
  DFFQX1 \desIn_r_reg[10]  ( .D(desIn[10]), .CK(n85), .Q(desIn_r[10]) );
  DFFQX1 \desIn_r_reg[8]  ( .D(desIn[8]), .CK(n85), .Q(desIn_r[8]) );
  DFFQX1 \desIn_r_reg[6]  ( .D(desIn[6]), .CK(n84), .Q(desIn_r[6]) );
  DFFQX1 \desIn_r_reg[4]  ( .D(desIn[4]), .CK(n84), .Q(desIn_r[4]) );
  DFFQX1 \desIn_r_reg[2]  ( .D(desIn[2]), .CK(n84), .Q(desIn_r[2]) );
  DFFQX1 \desIn_r_reg[0]  ( .D(desIn[0]), .CK(n84), .Q(desIn_r[0]) );
  DFFQX1 \L0_reg[1]  ( .D(desIn_r[7]), .CK(n84), .Q(L0[1]) );
  DFFQX1 \L0_reg[2]  ( .D(desIn_r[15]), .CK(n83), .Q(L0[2]) );
  DFFQX1 \L0_reg[3]  ( .D(desIn_r[23]), .CK(n83), .Q(L0[3]) );
  DFFQX1 \L0_reg[4]  ( .D(desIn_r[31]), .CK(n83), .Q(L0[4]) );
  DFFQX1 \L0_reg[5]  ( .D(desIn_r[39]), .CK(n83), .Q(L0[5]) );
  DFFQX1 \L0_reg[6]  ( .D(desIn_r[47]), .CK(n83), .Q(L0[6]) );
  DFFQX1 \L0_reg[7]  ( .D(desIn_r[55]), .CK(n83), .Q(L0[7]) );
  DFFQX1 \L0_reg[8]  ( .D(desIn_r[63]), .CK(n83), .Q(L0[8]) );
  DFFQX1 \L0_reg[9]  ( .D(desIn_r[5]), .CK(n83), .Q(L0[9]) );
  DFFQX1 \L0_reg[10]  ( .D(desIn_r[13]), .CK(n83), .Q(L0[10]) );
  DFFQX1 \L0_reg[11]  ( .D(desIn_r[21]), .CK(n82), .Q(L0[11]) );
  DFFQX1 \L0_reg[12]  ( .D(desIn_r[29]), .CK(n82), .Q(L0[12]) );
  DFFQX1 \L0_reg[13]  ( .D(desIn_r[37]), .CK(n82), .Q(L0[13]) );
  DFFQX1 \L0_reg[14]  ( .D(desIn_r[45]), .CK(n82), .Q(L0[14]) );
  DFFQX1 \L0_reg[15]  ( .D(desIn_r[53]), .CK(n82), .Q(L0[15]) );
  DFFQX1 \L0_reg[16]  ( .D(desIn_r[61]), .CK(n82), .Q(L0[16]) );
  DFFQX1 \L0_reg[17]  ( .D(desIn_r[3]), .CK(n82), .Q(L0[17]) );
  DFFQX1 \L0_reg[18]  ( .D(desIn_r[11]), .CK(n82), .Q(L0[18]) );
  DFFQX1 \L0_reg[19]  ( .D(desIn_r[19]), .CK(n82), .Q(L0[19]) );
  DFFQX1 \L0_reg[20]  ( .D(desIn_r[27]), .CK(n81), .Q(L0[20]) );
  DFFQX1 \L0_reg[21]  ( .D(desIn_r[35]), .CK(n81), .Q(L0[21]) );
  DFFQX1 \L0_reg[22]  ( .D(desIn_r[43]), .CK(n81), .Q(L0[22]) );
  DFFQX1 \L0_reg[23]  ( .D(desIn_r[51]), .CK(n81), .Q(L0[23]) );
  DFFQX1 \L0_reg[24]  ( .D(desIn_r[59]), .CK(n81), .Q(L0[24]) );
  DFFQX1 \L0_reg[25]  ( .D(desIn_r[1]), .CK(n81), .Q(L0[25]) );
  DFFQX1 \L0_reg[26]  ( .D(desIn_r[9]), .CK(n81), .Q(L0[26]) );
  DFFQX1 \L0_reg[27]  ( .D(desIn_r[17]), .CK(n81), .Q(L0[27]) );
  DFFQX1 \L0_reg[28]  ( .D(desIn_r[25]), .CK(n81), .Q(L0[28]) );
  DFFQX1 \L0_reg[29]  ( .D(desIn_r[33]), .CK(n80), .Q(L0[29]) );
  DFFQX1 \L0_reg[30]  ( .D(desIn_r[41]), .CK(n80), .Q(L0[30]) );
  DFFQX1 \L0_reg[31]  ( .D(desIn_r[49]), .CK(n80), .Q(L0[31]) );
  DFFQX1 \L0_reg[32]  ( .D(desIn_r[57]), .CK(n80), .Q(L0[32]) );
  DFFQX1 \L1_reg[1]  ( .D(R0[1]), .CK(n76), .Q(L1[1]) );
  DFFQX1 \L1_reg[2]  ( .D(R0[2]), .CK(n76), .Q(L1[2]) );
  DFFQX1 \L1_reg[3]  ( .D(R0[3]), .CK(n76), .Q(L1[3]) );
  DFFQX1 \L1_reg[4]  ( .D(R0[4]), .CK(n76), .Q(L1[4]) );
  DFFQX1 \L1_reg[5]  ( .D(R0[5]), .CK(n76), .Q(L1[5]) );
  DFFQX1 \L1_reg[6]  ( .D(R0[6]), .CK(n76), .Q(L1[6]) );
  DFFQX1 \L1_reg[7]  ( .D(R0[7]), .CK(n76), .Q(L1[7]) );
  DFFQX1 \L1_reg[8]  ( .D(R0[8]), .CK(n76), .Q(L1[8]) );
  DFFQX1 \L1_reg[9]  ( .D(R0[9]), .CK(n76), .Q(L1[9]) );
  DFFQX1 \L1_reg[10]  ( .D(R0[10]), .CK(n75), .Q(L1[10]) );
  DFFQX1 \L1_reg[11]  ( .D(R0[11]), .CK(n75), .Q(L1[11]) );
  DFFQX1 \L1_reg[12]  ( .D(R0[12]), .CK(n75), .Q(L1[12]) );
  DFFQX1 \L1_reg[13]  ( .D(R0[13]), .CK(n75), .Q(L1[13]) );
  DFFQX1 \L1_reg[14]  ( .D(R0[14]), .CK(n75), .Q(L1[14]) );
  DFFQX1 \L1_reg[15]  ( .D(R0[15]), .CK(n75), .Q(L1[15]) );
  DFFQX1 \L1_reg[16]  ( .D(R0[16]), .CK(n75), .Q(L1[16]) );
  DFFQX1 \L1_reg[17]  ( .D(R0[17]), .CK(n75), .Q(L1[17]) );
  DFFQX1 \L1_reg[18]  ( .D(R0[18]), .CK(n75), .Q(L1[18]) );
  DFFQX1 \L1_reg[19]  ( .D(R0[19]), .CK(n74), .Q(L1[19]) );
  DFFQX1 \L1_reg[20]  ( .D(R0[20]), .CK(n74), .Q(L1[20]) );
  DFFQX1 \L1_reg[21]  ( .D(R0[21]), .CK(n74), .Q(L1[21]) );
  DFFQX1 \L1_reg[22]  ( .D(R0[22]), .CK(n74), .Q(L1[22]) );
  DFFQX1 \L1_reg[23]  ( .D(R0[23]), .CK(n74), .Q(L1[23]) );
  DFFQX1 \L1_reg[24]  ( .D(R0[24]), .CK(n74), .Q(L1[24]) );
  DFFQX1 \L1_reg[25]  ( .D(R0[25]), .CK(n74), .Q(L1[25]) );
  DFFQX1 \L1_reg[26]  ( .D(R0[26]), .CK(n74), .Q(L1[26]) );
  DFFQX1 \L1_reg[27]  ( .D(R0[27]), .CK(n74), .Q(L1[27]) );
  DFFQX1 \L1_reg[28]  ( .D(R0[28]), .CK(n73), .Q(L1[28]) );
  DFFQX1 \L1_reg[29]  ( .D(R0[29]), .CK(n73), .Q(L1[29]) );
  DFFQX1 \L1_reg[30]  ( .D(R0[30]), .CK(n73), .Q(L1[30]) );
  DFFQX1 \L1_reg[31]  ( .D(R0[31]), .CK(n73), .Q(L1[31]) );
  DFFQX1 \L1_reg[32]  ( .D(R0[32]), .CK(n73), .Q(L1[32]) );
  DFFQX1 \L2_reg[1]  ( .D(R1[1]), .CK(n69), .Q(L2[1]) );
  DFFQX1 \L2_reg[2]  ( .D(R1[2]), .CK(n69), .Q(L2[2]) );
  DFFQX1 \L2_reg[3]  ( .D(R1[3]), .CK(n69), .Q(L2[3]) );
  DFFQX1 \L2_reg[4]  ( .D(R1[4]), .CK(n69), .Q(L2[4]) );
  DFFQX1 \L2_reg[5]  ( .D(R1[5]), .CK(n69), .Q(L2[5]) );
  DFFQX1 \L2_reg[6]  ( .D(R1[6]), .CK(n69), .Q(L2[6]) );
  DFFQX1 \L2_reg[7]  ( .D(R1[7]), .CK(n69), .Q(L2[7]) );
  DFFQX1 \L2_reg[8]  ( .D(R1[8]), .CK(n69), .Q(L2[8]) );
  DFFQX1 \L2_reg[9]  ( .D(R1[9]), .CK(n68), .Q(L2[9]) );
  DFFQX1 \L2_reg[10]  ( .D(R1[10]), .CK(n68), .Q(L2[10]) );
  DFFQX1 \L2_reg[11]  ( .D(R1[11]), .CK(n68), .Q(L2[11]) );
  DFFQX1 \L2_reg[12]  ( .D(R1[12]), .CK(n68), .Q(L2[12]) );
  DFFQX1 \L2_reg[13]  ( .D(R1[13]), .CK(n68), .Q(L2[13]) );
  DFFQX1 \L2_reg[14]  ( .D(R1[14]), .CK(n68), .Q(L2[14]) );
  DFFQX1 \L2_reg[15]  ( .D(R1[15]), .CK(n68), .Q(L2[15]) );
  DFFQX1 \L2_reg[16]  ( .D(R1[16]), .CK(n68), .Q(L2[16]) );
  DFFQX1 \L2_reg[17]  ( .D(R1[17]), .CK(n68), .Q(L2[17]) );
  DFFQX1 \L2_reg[18]  ( .D(R1[18]), .CK(n67), .Q(L2[18]) );
  DFFQX1 \L2_reg[19]  ( .D(R1[19]), .CK(n67), .Q(L2[19]) );
  DFFQX1 \L2_reg[20]  ( .D(R1[20]), .CK(n67), .Q(L2[20]) );
  DFFQX1 \L2_reg[21]  ( .D(R1[21]), .CK(n67), .Q(L2[21]) );
  DFFQX1 \L2_reg[22]  ( .D(R1[22]), .CK(n67), .Q(L2[22]) );
  DFFQX1 \L2_reg[23]  ( .D(R1[23]), .CK(n67), .Q(L2[23]) );
  DFFQX1 \L2_reg[24]  ( .D(R1[24]), .CK(n67), .Q(L2[24]) );
  DFFQX1 \L2_reg[25]  ( .D(R1[25]), .CK(n67), .Q(L2[25]) );
  DFFQX1 \L2_reg[26]  ( .D(R1[26]), .CK(n67), .Q(L2[26]) );
  DFFQX1 \L2_reg[27]  ( .D(R1[27]), .CK(n66), .Q(L2[27]) );
  DFFQX1 \L2_reg[28]  ( .D(R1[28]), .CK(n66), .Q(L2[28]) );
  DFFQX1 \L2_reg[29]  ( .D(R1[29]), .CK(n66), .Q(L2[29]) );
  DFFQX1 \L2_reg[30]  ( .D(R1[30]), .CK(n66), .Q(L2[30]) );
  DFFQX1 \L2_reg[31]  ( .D(R1[31]), .CK(n66), .Q(L2[31]) );
  DFFQX1 \L2_reg[32]  ( .D(R1[32]), .CK(n66), .Q(L2[32]) );
  DFFQX1 \L3_reg[1]  ( .D(R2[1]), .CK(n62), .Q(L3[1]) );
  DFFQX1 \L3_reg[2]  ( .D(R2[2]), .CK(n62), .Q(L3[2]) );
  DFFQX1 \L3_reg[3]  ( .D(R2[3]), .CK(n62), .Q(L3[3]) );
  DFFQX1 \L3_reg[4]  ( .D(R2[4]), .CK(n62), .Q(L3[4]) );
  DFFQX1 \L3_reg[5]  ( .D(R2[5]), .CK(n62), .Q(L3[5]) );
  DFFQX1 \L3_reg[6]  ( .D(R2[6]), .CK(n62), .Q(L3[6]) );
  DFFQX1 \L3_reg[7]  ( .D(R2[7]), .CK(n62), .Q(L3[7]) );
  DFFQX1 \L3_reg[8]  ( .D(R2[8]), .CK(n61), .Q(L3[8]) );
  DFFQX1 \L3_reg[9]  ( .D(R2[9]), .CK(n61), .Q(L3[9]) );
  DFFQX1 \L3_reg[10]  ( .D(R2[10]), .CK(n61), .Q(L3[10]) );
  DFFQX1 \L3_reg[11]  ( .D(R2[11]), .CK(n61), .Q(L3[11]) );
  DFFQX1 \L3_reg[12]  ( .D(R2[12]), .CK(n61), .Q(L3[12]) );
  DFFQX1 \L3_reg[13]  ( .D(R2[13]), .CK(n61), .Q(L3[13]) );
  DFFQX1 \L3_reg[14]  ( .D(R2[14]), .CK(n61), .Q(L3[14]) );
  DFFQX1 \L3_reg[15]  ( .D(R2[15]), .CK(n61), .Q(L3[15]) );
  DFFQX1 \L3_reg[16]  ( .D(R2[16]), .CK(n61), .Q(L3[16]) );
  DFFQX1 \L3_reg[17]  ( .D(R2[17]), .CK(n60), .Q(L3[17]) );
  DFFQX1 \L3_reg[18]  ( .D(R2[18]), .CK(n60), .Q(L3[18]) );
  DFFQX1 \L3_reg[19]  ( .D(R2[19]), .CK(n60), .Q(L3[19]) );
  DFFQX1 \L3_reg[20]  ( .D(R2[20]), .CK(n60), .Q(L3[20]) );
  DFFQX1 \L3_reg[21]  ( .D(R2[21]), .CK(n60), .Q(L3[21]) );
  DFFQX1 \L3_reg[22]  ( .D(R2[22]), .CK(n60), .Q(L3[22]) );
  DFFQX1 \L3_reg[23]  ( .D(R2[23]), .CK(n60), .Q(L3[23]) );
  DFFQX1 \L3_reg[24]  ( .D(R2[24]), .CK(n60), .Q(L3[24]) );
  DFFQX1 \L3_reg[25]  ( .D(R2[25]), .CK(n60), .Q(L3[25]) );
  DFFQX1 \L3_reg[26]  ( .D(R2[26]), .CK(n59), .Q(L3[26]) );
  DFFQX1 \L3_reg[27]  ( .D(R2[27]), .CK(n59), .Q(L3[27]) );
  DFFQX1 \L3_reg[28]  ( .D(R2[28]), .CK(n59), .Q(L3[28]) );
  DFFQX1 \L3_reg[29]  ( .D(R2[29]), .CK(n59), .Q(L3[29]) );
  DFFQX1 \L3_reg[30]  ( .D(R2[30]), .CK(n59), .Q(L3[30]) );
  DFFQX1 \L3_reg[31]  ( .D(R2[31]), .CK(n59), .Q(L3[31]) );
  DFFQX1 \L3_reg[32]  ( .D(R2[32]), .CK(n59), .Q(L3[32]) );
  DFFQX1 \L4_reg[1]  ( .D(R3[1]), .CK(n55), .Q(L4[1]) );
  DFFQX1 \L4_reg[2]  ( .D(R3[2]), .CK(n55), .Q(L4[2]) );
  DFFQX1 \L4_reg[3]  ( .D(R3[3]), .CK(n55), .Q(L4[3]) );
  DFFQX1 \L4_reg[4]  ( .D(R3[4]), .CK(n55), .Q(L4[4]) );
  DFFQX1 \L4_reg[5]  ( .D(R3[5]), .CK(n55), .Q(L4[5]) );
  DFFQX1 \L4_reg[6]  ( .D(R3[6]), .CK(n55), .Q(L4[6]) );
  DFFQX1 \L4_reg[7]  ( .D(R3[7]), .CK(n54), .Q(L4[7]) );
  DFFQX1 \L4_reg[8]  ( .D(R3[8]), .CK(n54), .Q(L4[8]) );
  DFFQX1 \L4_reg[9]  ( .D(R3[9]), .CK(n54), .Q(L4[9]) );
  DFFQX1 \L4_reg[10]  ( .D(R3[10]), .CK(n54), .Q(L4[10]) );
  DFFQX1 \L4_reg[11]  ( .D(R3[11]), .CK(n54), .Q(L4[11]) );
  DFFQX1 \L4_reg[12]  ( .D(R3[12]), .CK(n54), .Q(L4[12]) );
  DFFQX1 \L4_reg[13]  ( .D(R3[13]), .CK(n54), .Q(L4[13]) );
  DFFQX1 \L4_reg[14]  ( .D(R3[14]), .CK(n54), .Q(L4[14]) );
  DFFQX1 \L4_reg[15]  ( .D(R3[15]), .CK(n54), .Q(L4[15]) );
  DFFQX1 \L4_reg[16]  ( .D(R3[16]), .CK(n53), .Q(L4[16]) );
  DFFQX1 \L4_reg[17]  ( .D(R3[17]), .CK(n53), .Q(L4[17]) );
  DFFQX1 \L4_reg[18]  ( .D(R3[18]), .CK(n53), .Q(L4[18]) );
  DFFQX1 \L4_reg[19]  ( .D(R3[19]), .CK(n53), .Q(L4[19]) );
  DFFQX1 \L4_reg[20]  ( .D(R3[20]), .CK(n53), .Q(L4[20]) );
  DFFQX1 \L4_reg[21]  ( .D(R3[21]), .CK(n53), .Q(L4[21]) );
  DFFQX1 \L4_reg[22]  ( .D(R3[22]), .CK(n53), .Q(L4[22]) );
  DFFQX1 \L4_reg[23]  ( .D(R3[23]), .CK(n53), .Q(L4[23]) );
  DFFQX1 \L4_reg[24]  ( .D(R3[24]), .CK(n53), .Q(L4[24]) );
  DFFQX1 \L4_reg[25]  ( .D(R3[25]), .CK(n52), .Q(L4[25]) );
  DFFQX1 \L4_reg[26]  ( .D(R3[26]), .CK(n52), .Q(L4[26]) );
  DFFQX1 \L4_reg[27]  ( .D(R3[27]), .CK(n52), .Q(L4[27]) );
  DFFQX1 \L4_reg[28]  ( .D(R3[28]), .CK(n52), .Q(L4[28]) );
  DFFQX1 \L4_reg[29]  ( .D(R3[29]), .CK(n52), .Q(L4[29]) );
  DFFQX1 \L4_reg[30]  ( .D(R3[30]), .CK(n52), .Q(L4[30]) );
  DFFQX1 \L4_reg[31]  ( .D(R3[31]), .CK(n52), .Q(L4[31]) );
  DFFQX1 \L4_reg[32]  ( .D(R3[32]), .CK(n52), .Q(L4[32]) );
  DFFQX1 \L5_reg[1]  ( .D(R4[1]), .CK(n48), .Q(L5[1]) );
  DFFQX1 \L5_reg[2]  ( .D(R4[2]), .CK(n48), .Q(L5[2]) );
  DFFQX1 \L5_reg[3]  ( .D(R4[3]), .CK(n48), .Q(L5[3]) );
  DFFQX1 \L5_reg[4]  ( .D(R4[4]), .CK(n48), .Q(L5[4]) );
  DFFQX1 \L5_reg[5]  ( .D(R4[5]), .CK(n48), .Q(L5[5]) );
  DFFQX1 \L5_reg[6]  ( .D(R4[6]), .CK(n47), .Q(L5[6]) );
  DFFQX1 \L5_reg[7]  ( .D(R4[7]), .CK(n47), .Q(L5[7]) );
  DFFQX1 \L5_reg[8]  ( .D(R4[8]), .CK(n47), .Q(L5[8]) );
  DFFQX1 \L5_reg[9]  ( .D(R4[9]), .CK(n47), .Q(L5[9]) );
  DFFQX1 \L5_reg[10]  ( .D(R4[10]), .CK(n47), .Q(L5[10]) );
  DFFQX1 \L5_reg[11]  ( .D(R4[11]), .CK(n47), .Q(L5[11]) );
  DFFQX1 \L5_reg[12]  ( .D(R4[12]), .CK(n47), .Q(L5[12]) );
  DFFQX1 \L5_reg[13]  ( .D(R4[13]), .CK(n47), .Q(L5[13]) );
  DFFQX1 \L5_reg[14]  ( .D(R4[14]), .CK(n47), .Q(L5[14]) );
  DFFQX1 \L5_reg[15]  ( .D(R4[15]), .CK(n46), .Q(L5[15]) );
  DFFQX1 \L5_reg[16]  ( .D(R4[16]), .CK(n46), .Q(L5[16]) );
  DFFQX1 \L5_reg[17]  ( .D(R4[17]), .CK(n46), .Q(L5[17]) );
  DFFQX1 \L5_reg[18]  ( .D(R4[18]), .CK(n46), .Q(L5[18]) );
  DFFQX1 \L5_reg[19]  ( .D(R4[19]), .CK(n46), .Q(L5[19]) );
  DFFQX1 \L5_reg[20]  ( .D(R4[20]), .CK(n46), .Q(L5[20]) );
  DFFQX1 \L5_reg[21]  ( .D(R4[21]), .CK(n46), .Q(L5[21]) );
  DFFQX1 \L5_reg[22]  ( .D(R4[22]), .CK(n46), .Q(L5[22]) );
  DFFQX1 \L5_reg[23]  ( .D(R4[23]), .CK(n46), .Q(L5[23]) );
  DFFQX1 \L5_reg[24]  ( .D(R4[24]), .CK(n45), .Q(L5[24]) );
  DFFQX1 \L5_reg[25]  ( .D(R4[25]), .CK(n45), .Q(L5[25]) );
  DFFQX1 \L5_reg[26]  ( .D(R4[26]), .CK(n45), .Q(L5[26]) );
  DFFQX1 \L5_reg[27]  ( .D(R4[27]), .CK(n45), .Q(L5[27]) );
  DFFQX1 \L5_reg[28]  ( .D(R4[28]), .CK(n45), .Q(L5[28]) );
  DFFQX1 \L5_reg[29]  ( .D(R4[29]), .CK(n45), .Q(L5[29]) );
  DFFQX1 \L5_reg[30]  ( .D(R4[30]), .CK(n45), .Q(L5[30]) );
  DFFQX1 \L5_reg[31]  ( .D(R4[31]), .CK(n45), .Q(L5[31]) );
  DFFQX1 \L5_reg[32]  ( .D(R4[32]), .CK(n45), .Q(L5[32]) );
  DFFQX1 \L6_reg[1]  ( .D(R5[1]), .CK(n41), .Q(L6[1]) );
  DFFQX1 \L6_reg[2]  ( .D(R5[2]), .CK(n41), .Q(L6[2]) );
  DFFQX1 \L6_reg[3]  ( .D(R5[3]), .CK(n41), .Q(L6[3]) );
  DFFQX1 \L6_reg[4]  ( .D(R5[4]), .CK(n41), .Q(L6[4]) );
  DFFQX1 \L6_reg[5]  ( .D(R5[5]), .CK(n40), .Q(L6[5]) );
  DFFQX1 \L6_reg[6]  ( .D(R5[6]), .CK(n40), .Q(L6[6]) );
  DFFQX1 \L6_reg[7]  ( .D(R5[7]), .CK(n40), .Q(L6[7]) );
  DFFQX1 \L6_reg[8]  ( .D(R5[8]), .CK(n40), .Q(L6[8]) );
  DFFQX1 \L6_reg[9]  ( .D(R5[9]), .CK(n40), .Q(L6[9]) );
  DFFQX1 \L6_reg[10]  ( .D(R5[10]), .CK(n40), .Q(L6[10]) );
  DFFQX1 \L6_reg[11]  ( .D(R5[11]), .CK(n40), .Q(L6[11]) );
  DFFQX1 \L6_reg[12]  ( .D(R5[12]), .CK(n40), .Q(L6[12]) );
  DFFQX1 \L6_reg[13]  ( .D(R5[13]), .CK(n40), .Q(L6[13]) );
  DFFQX1 \L6_reg[14]  ( .D(R5[14]), .CK(n39), .Q(L6[14]) );
  DFFQX1 \L6_reg[15]  ( .D(R5[15]), .CK(n39), .Q(L6[15]) );
  DFFQX1 \L6_reg[16]  ( .D(R5[16]), .CK(n39), .Q(L6[16]) );
  DFFQX1 \L6_reg[17]  ( .D(R5[17]), .CK(n39), .Q(L6[17]) );
  DFFQX1 \L6_reg[18]  ( .D(R5[18]), .CK(n39), .Q(L6[18]) );
  DFFQX1 \L6_reg[19]  ( .D(R5[19]), .CK(n39), .Q(L6[19]) );
  DFFQX1 \L6_reg[20]  ( .D(R5[20]), .CK(n39), .Q(L6[20]) );
  DFFQX1 \L6_reg[21]  ( .D(R5[21]), .CK(n39), .Q(L6[21]) );
  DFFQX1 \L6_reg[22]  ( .D(R5[22]), .CK(n39), .Q(L6[22]) );
  DFFQX1 \L6_reg[23]  ( .D(R5[23]), .CK(n38), .Q(L6[23]) );
  DFFQX1 \L6_reg[24]  ( .D(R5[24]), .CK(n38), .Q(L6[24]) );
  DFFQX1 \L6_reg[25]  ( .D(R5[25]), .CK(n38), .Q(L6[25]) );
  DFFQX1 \L6_reg[26]  ( .D(R5[26]), .CK(n38), .Q(L6[26]) );
  DFFQX1 \L6_reg[27]  ( .D(R5[27]), .CK(n38), .Q(L6[27]) );
  DFFQX1 \L6_reg[28]  ( .D(R5[28]), .CK(n38), .Q(L6[28]) );
  DFFQX1 \L6_reg[29]  ( .D(R5[29]), .CK(n38), .Q(L6[29]) );
  DFFQX1 \L6_reg[30]  ( .D(R5[30]), .CK(n38), .Q(L6[30]) );
  DFFQX1 \L6_reg[31]  ( .D(R5[31]), .CK(n38), .Q(L6[31]) );
  DFFQX1 \L6_reg[32]  ( .D(R5[32]), .CK(n37), .Q(L6[32]) );
  DFFQX1 \L7_reg[1]  ( .D(R6[1]), .CK(n34), .Q(L7[1]) );
  DFFQX1 \L7_reg[2]  ( .D(R6[2]), .CK(n34), .Q(L7[2]) );
  DFFQX1 \L7_reg[3]  ( .D(R6[3]), .CK(n34), .Q(L7[3]) );
  DFFQX1 \L7_reg[4]  ( .D(R6[4]), .CK(n33), .Q(L7[4]) );
  DFFQX1 \L7_reg[5]  ( .D(R6[5]), .CK(n33), .Q(L7[5]) );
  DFFQX1 \L7_reg[6]  ( .D(R6[6]), .CK(n33), .Q(L7[6]) );
  DFFQX1 \L7_reg[7]  ( .D(R6[7]), .CK(n33), .Q(L7[7]) );
  DFFQX1 \L7_reg[8]  ( .D(R6[8]), .CK(n33), .Q(L7[8]) );
  DFFQX1 \L7_reg[9]  ( .D(R6[9]), .CK(n33), .Q(L7[9]) );
  DFFQX1 \L7_reg[10]  ( .D(R6[10]), .CK(n33), .Q(L7[10]) );
  DFFQX1 \L7_reg[11]  ( .D(R6[11]), .CK(n33), .Q(L7[11]) );
  DFFQX1 \L7_reg[12]  ( .D(R6[12]), .CK(n33), .Q(L7[12]) );
  DFFQX1 \L7_reg[13]  ( .D(R6[13]), .CK(n32), .Q(L7[13]) );
  DFFQX1 \L7_reg[14]  ( .D(R6[14]), .CK(n32), .Q(L7[14]) );
  DFFQX1 \L7_reg[15]  ( .D(R6[15]), .CK(n32), .Q(L7[15]) );
  DFFQX1 \L7_reg[16]  ( .D(R6[16]), .CK(n32), .Q(L7[16]) );
  DFFQX1 \L7_reg[17]  ( .D(R6[17]), .CK(n32), .Q(L7[17]) );
  DFFQX1 \L7_reg[18]  ( .D(R6[18]), .CK(n32), .Q(L7[18]) );
  DFFQX1 \L7_reg[19]  ( .D(R6[19]), .CK(n32), .Q(L7[19]) );
  DFFQX1 \L7_reg[20]  ( .D(R6[20]), .CK(n32), .Q(L7[20]) );
  DFFQX1 \L7_reg[21]  ( .D(R6[21]), .CK(n32), .Q(L7[21]) );
  DFFQX1 \L7_reg[22]  ( .D(R6[22]), .CK(n31), .Q(L7[22]) );
  DFFQX1 \L7_reg[23]  ( .D(R6[23]), .CK(n31), .Q(L7[23]) );
  DFFQX1 \L7_reg[24]  ( .D(R6[24]), .CK(n31), .Q(L7[24]) );
  DFFQX1 \L7_reg[25]  ( .D(R6[25]), .CK(n31), .Q(L7[25]) );
  DFFQX1 \L7_reg[26]  ( .D(R6[26]), .CK(n31), .Q(L7[26]) );
  DFFQX1 \L7_reg[27]  ( .D(R6[27]), .CK(n31), .Q(L7[27]) );
  DFFQX1 \L7_reg[28]  ( .D(R6[28]), .CK(n31), .Q(L7[28]) );
  DFFQX1 \L7_reg[29]  ( .D(R6[29]), .CK(n31), .Q(L7[29]) );
  DFFQX1 \L7_reg[30]  ( .D(R6[30]), .CK(n31), .Q(L7[30]) );
  DFFQX1 \L7_reg[31]  ( .D(R6[31]), .CK(n30), .Q(L7[31]) );
  DFFQX1 \L7_reg[32]  ( .D(R6[32]), .CK(n30), .Q(L7[32]) );
  DFFQX1 \L8_reg[1]  ( .D(R7[1]), .CK(n27), .Q(L8[1]) );
  DFFQX1 \L8_reg[2]  ( .D(R7[2]), .CK(n27), .Q(L8[2]) );
  DFFQX1 \L8_reg[3]  ( .D(R7[3]), .CK(n26), .Q(L8[3]) );
  DFFQX1 \L8_reg[4]  ( .D(R7[4]), .CK(n26), .Q(L8[4]) );
  DFFQX1 \L8_reg[5]  ( .D(R7[5]), .CK(n26), .Q(L8[5]) );
  DFFQX1 \L8_reg[6]  ( .D(R7[6]), .CK(n26), .Q(L8[6]) );
  DFFQX1 \L8_reg[7]  ( .D(R7[7]), .CK(n26), .Q(L8[7]) );
  DFFQX1 \L8_reg[8]  ( .D(R7[8]), .CK(n26), .Q(L8[8]) );
  DFFQX1 \L8_reg[9]  ( .D(R7[9]), .CK(n26), .Q(L8[9]) );
  DFFQX1 \L8_reg[10]  ( .D(R7[10]), .CK(n26), .Q(L8[10]) );
  DFFQX1 \L8_reg[11]  ( .D(R7[11]), .CK(n26), .Q(L8[11]) );
  DFFQX1 \L8_reg[12]  ( .D(R7[12]), .CK(n25), .Q(L8[12]) );
  DFFQX1 \L8_reg[13]  ( .D(R7[13]), .CK(n25), .Q(L8[13]) );
  DFFQX1 \L8_reg[14]  ( .D(R7[14]), .CK(n25), .Q(L8[14]) );
  DFFQX1 \L8_reg[15]  ( .D(R7[15]), .CK(n25), .Q(L8[15]) );
  DFFQX1 \L8_reg[16]  ( .D(R7[16]), .CK(n25), .Q(L8[16]) );
  DFFQX1 \L8_reg[17]  ( .D(R7[17]), .CK(n25), .Q(L8[17]) );
  DFFQX1 \L8_reg[18]  ( .D(R7[18]), .CK(n25), .Q(L8[18]) );
  DFFQX1 \L8_reg[19]  ( .D(R7[19]), .CK(n25), .Q(L8[19]) );
  DFFQX1 \L8_reg[20]  ( .D(R7[20]), .CK(n25), .Q(L8[20]) );
  DFFQX1 \L8_reg[21]  ( .D(R7[21]), .CK(n24), .Q(L8[21]) );
  DFFQX1 \L8_reg[22]  ( .D(R7[22]), .CK(n24), .Q(L8[22]) );
  DFFQX1 \L8_reg[23]  ( .D(R7[23]), .CK(n24), .Q(L8[23]) );
  DFFQX1 \L8_reg[24]  ( .D(R7[24]), .CK(n24), .Q(L8[24]) );
  DFFQX1 \L8_reg[25]  ( .D(R7[25]), .CK(n24), .Q(L8[25]) );
  DFFQX1 \L8_reg[26]  ( .D(R7[26]), .CK(n24), .Q(L8[26]) );
  DFFQX1 \L8_reg[27]  ( .D(R7[27]), .CK(n24), .Q(L8[27]) );
  DFFQX1 \L8_reg[28]  ( .D(R7[28]), .CK(n24), .Q(L8[28]) );
  DFFQX1 \L8_reg[29]  ( .D(R7[29]), .CK(n24), .Q(L8[29]) );
  DFFQX1 \L8_reg[30]  ( .D(R7[30]), .CK(n23), .Q(L8[30]) );
  DFFQX1 \L8_reg[31]  ( .D(R7[31]), .CK(n23), .Q(L8[31]) );
  DFFQX1 \L8_reg[32]  ( .D(R7[32]), .CK(n23), .Q(L8[32]) );
  DFFQX1 \L9_reg[1]  ( .D(R8[1]), .CK(n20), .Q(L9[1]) );
  DFFQX1 \L9_reg[2]  ( .D(R8[2]), .CK(n19), .Q(L9[2]) );
  DFFQX1 \L9_reg[3]  ( .D(R8[3]), .CK(n19), .Q(L9[3]) );
  DFFQX1 \L9_reg[4]  ( .D(R8[4]), .CK(n19), .Q(L9[4]) );
  DFFQX1 \L9_reg[5]  ( .D(R8[5]), .CK(n19), .Q(L9[5]) );
  DFFQX1 \L9_reg[6]  ( .D(R8[6]), .CK(n19), .Q(L9[6]) );
  DFFQX1 \L9_reg[7]  ( .D(R8[7]), .CK(n19), .Q(L9[7]) );
  DFFQX1 \L9_reg[8]  ( .D(R8[8]), .CK(n19), .Q(L9[8]) );
  DFFQX1 \L9_reg[9]  ( .D(R8[9]), .CK(n19), .Q(L9[9]) );
  DFFQX1 \L9_reg[10]  ( .D(R8[10]), .CK(n19), .Q(L9[10]) );
  DFFQX1 \L9_reg[11]  ( .D(R8[11]), .CK(n18), .Q(L9[11]) );
  DFFQX1 \L9_reg[12]  ( .D(R8[12]), .CK(n18), .Q(L9[12]) );
  DFFQX1 \L9_reg[13]  ( .D(R8[13]), .CK(n18), .Q(L9[13]) );
  DFFQX1 \L9_reg[14]  ( .D(R8[14]), .CK(n18), .Q(L9[14]) );
  DFFQX1 \L9_reg[15]  ( .D(R8[15]), .CK(n18), .Q(L9[15]) );
  DFFQX1 \L9_reg[16]  ( .D(R8[16]), .CK(n18), .Q(L9[16]) );
  DFFQX1 \L9_reg[17]  ( .D(R8[17]), .CK(n18), .Q(L9[17]) );
  DFFQX1 \L9_reg[18]  ( .D(R8[18]), .CK(n18), .Q(L9[18]) );
  DFFQX1 \L9_reg[19]  ( .D(R8[19]), .CK(n18), .Q(L9[19]) );
  DFFQX1 \L9_reg[20]  ( .D(R8[20]), .CK(n17), .Q(L9[20]) );
  DFFQX1 \L9_reg[21]  ( .D(R8[21]), .CK(n17), .Q(L9[21]) );
  DFFQX1 \L9_reg[22]  ( .D(R8[22]), .CK(n17), .Q(L9[22]) );
  DFFQX1 \L9_reg[23]  ( .D(R8[23]), .CK(n17), .Q(L9[23]) );
  DFFQX1 \L9_reg[24]  ( .D(R8[24]), .CK(n17), .Q(L9[24]) );
  DFFQX1 \L9_reg[25]  ( .D(R8[25]), .CK(n17), .Q(L9[25]) );
  DFFQX1 \L9_reg[26]  ( .D(R8[26]), .CK(n17), .Q(L9[26]) );
  DFFQX1 \L9_reg[27]  ( .D(R8[27]), .CK(n17), .Q(L9[27]) );
  DFFQX1 \L9_reg[28]  ( .D(R8[28]), .CK(n17), .Q(L9[28]) );
  DFFQX1 \L9_reg[29]  ( .D(R8[29]), .CK(n16), .Q(L9[29]) );
  DFFQX1 \L9_reg[30]  ( .D(R8[30]), .CK(n16), .Q(L9[30]) );
  DFFQX1 \L9_reg[31]  ( .D(R8[31]), .CK(n16), .Q(L9[31]) );
  DFFQX1 \L9_reg[32]  ( .D(R8[32]), .CK(n16), .Q(L9[32]) );
  DFFQX1 \L10_reg[1]  ( .D(R9[1]), .CK(n12), .Q(L10[1]) );
  DFFQX1 \L10_reg[2]  ( .D(R9[2]), .CK(n12), .Q(L10[2]) );
  DFFQX1 \L10_reg[3]  ( .D(R9[3]), .CK(n12), .Q(L10[3]) );
  DFFQX1 \L10_reg[4]  ( .D(R9[4]), .CK(n12), .Q(L10[4]) );
  DFFQX1 \L10_reg[5]  ( .D(R9[5]), .CK(n12), .Q(L10[5]) );
  DFFQX1 \L10_reg[6]  ( .D(R9[6]), .CK(n12), .Q(L10[6]) );
  DFFQX1 \L10_reg[7]  ( .D(R9[7]), .CK(n12), .Q(L10[7]) );
  DFFQX1 \L10_reg[8]  ( .D(R9[8]), .CK(n12), .Q(L10[8]) );
  DFFQX1 \L10_reg[9]  ( .D(R9[9]), .CK(n12), .Q(L10[9]) );
  DFFQX1 \L10_reg[10]  ( .D(R9[10]), .CK(n11), .Q(L10[10]) );
  DFFQX1 \L10_reg[11]  ( .D(R9[11]), .CK(n11), .Q(L10[11]) );
  DFFQX1 \L10_reg[12]  ( .D(R9[12]), .CK(n11), .Q(L10[12]) );
  DFFQX1 \L10_reg[13]  ( .D(R9[13]), .CK(n11), .Q(L10[13]) );
  DFFQX1 \L10_reg[14]  ( .D(R9[14]), .CK(n11), .Q(L10[14]) );
  DFFQX1 \L10_reg[15]  ( .D(R9[15]), .CK(n11), .Q(L10[15]) );
  DFFQX1 \L10_reg[16]  ( .D(R9[16]), .CK(n11), .Q(L10[16]) );
  DFFQX1 \L10_reg[17]  ( .D(R9[17]), .CK(n11), .Q(L10[17]) );
  DFFQX1 \L10_reg[18]  ( .D(R9[18]), .CK(n11), .Q(L10[18]) );
  DFFQX1 \L10_reg[19]  ( .D(R9[19]), .CK(n10), .Q(L10[19]) );
  DFFQX1 \L10_reg[20]  ( .D(R9[20]), .CK(n10), .Q(L10[20]) );
  DFFQX1 \L10_reg[21]  ( .D(R9[21]), .CK(n10), .Q(L10[21]) );
  DFFQX1 \L10_reg[22]  ( .D(R9[22]), .CK(n10), .Q(L10[22]) );
  DFFQX1 \L10_reg[23]  ( .D(R9[23]), .CK(n10), .Q(L10[23]) );
  DFFQX1 \L10_reg[24]  ( .D(R9[24]), .CK(n10), .Q(L10[24]) );
  DFFQX1 \L10_reg[25]  ( .D(R9[25]), .CK(n10), .Q(L10[25]) );
  DFFQX1 \L10_reg[26]  ( .D(R9[26]), .CK(n10), .Q(L10[26]) );
  DFFQX1 \L10_reg[27]  ( .D(R9[27]), .CK(n10), .Q(L10[27]) );
  DFFQX1 \L10_reg[28]  ( .D(R9[28]), .CK(n9), .Q(L10[28]) );
  DFFQX1 \L10_reg[29]  ( .D(R9[29]), .CK(n9), .Q(L10[29]) );
  DFFQX1 \L10_reg[30]  ( .D(R9[30]), .CK(n9), .Q(L10[30]) );
  DFFQX1 \L10_reg[31]  ( .D(R9[31]), .CK(n9), .Q(L10[31]) );
  DFFQX1 \L10_reg[32]  ( .D(R9[32]), .CK(n9), .Q(L10[32]) );
  DFFQX1 \L11_reg[1]  ( .D(R10[1]), .CK(n5), .Q(L11[1]) );
  DFFQX1 \L11_reg[2]  ( .D(R10[2]), .CK(n5), .Q(L11[2]) );
  DFFQX1 \L11_reg[3]  ( .D(R10[3]), .CK(n5), .Q(L11[3]) );
  DFFQX1 \L11_reg[4]  ( .D(R10[4]), .CK(n5), .Q(L11[4]) );
  DFFQX1 \L11_reg[5]  ( .D(R10[5]), .CK(n5), .Q(L11[5]) );
  DFFQX1 \L11_reg[6]  ( .D(R10[6]), .CK(n5), .Q(L11[6]) );
  DFFQX1 \L11_reg[7]  ( .D(R10[7]), .CK(n5), .Q(L11[7]) );
  DFFQX1 \L11_reg[8]  ( .D(R10[8]), .CK(n5), .Q(L11[8]) );
  DFFQX1 \L11_reg[9]  ( .D(R10[9]), .CK(n4), .Q(L11[9]) );
  DFFQX1 \L11_reg[10]  ( .D(R10[10]), .CK(n4), .Q(L11[10]) );
  DFFQX1 \L11_reg[11]  ( .D(R10[11]), .CK(n4), .Q(L11[11]) );
  DFFQX1 \L11_reg[12]  ( .D(R10[12]), .CK(n4), .Q(L11[12]) );
  DFFQX1 \L11_reg[13]  ( .D(R10[13]), .CK(n4), .Q(L11[13]) );
  DFFQX1 \L11_reg[14]  ( .D(R10[14]), .CK(n4), .Q(L11[14]) );
  DFFQX1 \L11_reg[15]  ( .D(R10[15]), .CK(n4), .Q(L11[15]) );
  DFFQX1 \L11_reg[16]  ( .D(R10[16]), .CK(n4), .Q(L11[16]) );
  DFFQX1 \L11_reg[17]  ( .D(R10[17]), .CK(n4), .Q(L11[17]) );
  DFFQX1 \L11_reg[18]  ( .D(R10[18]), .CK(n90), .Q(L11[18]) );
  DFFQX1 \L11_reg[19]  ( .D(R10[19]), .CK(n20), .Q(L11[19]) );
  DFFQX1 \L11_reg[20]  ( .D(R10[20]), .CK(n13), .Q(L11[20]) );
  DFFQX1 \L11_reg[21]  ( .D(R10[21]), .CK(n6), .Q(L11[21]) );
  DFFQX1 \L11_reg[22]  ( .D(R10[22]), .CK(n77), .Q(L11[22]) );
  DFFQX1 \L11_reg[23]  ( .D(R10[23]), .CK(n70), .Q(L11[23]) );
  DFFQX1 \L11_reg[24]  ( .D(R10[24]), .CK(n63), .Q(L11[24]) );
  DFFQX1 \L11_reg[25]  ( .D(R10[25]), .CK(n58), .Q(L11[25]) );
  DFFQX1 \L11_reg[26]  ( .D(R10[26]), .CK(n56), .Q(L11[26]) );
  DFFQX1 \L11_reg[27]  ( .D(R10[27]), .CK(n72), .Q(L11[27]) );
  DFFQX1 \L11_reg[28]  ( .D(R10[28]), .CK(n71), .Q(L11[28]) );
  DFFQX1 \L11_reg[29]  ( .D(R10[29]), .CK(n65), .Q(L11[29]) );
  DFFQX1 \L11_reg[30]  ( .D(R10[30]), .CK(n64), .Q(L11[30]) );
  DFFQX1 \L11_reg[31]  ( .D(R10[31]), .CK(n50), .Q(L11[31]) );
  DFFQX1 \L11_reg[32]  ( .D(R10[32]), .CK(n43), .Q(L11[32]) );
  DFFQX1 \L12_reg[1]  ( .D(R11[1]), .CK(n67), .Q(L12[1]) );
  DFFQX1 \L12_reg[2]  ( .D(R11[2]), .CK(n66), .Q(L12[2]) );
  DFFQX1 \L12_reg[3]  ( .D(R11[3]), .CK(n62), .Q(L12[3]) );
  DFFQX1 \L12_reg[4]  ( .D(R11[4]), .CK(n61), .Q(L12[4]) );
  DFFQX1 \L12_reg[5]  ( .D(R11[5]), .CK(n60), .Q(L12[5]) );
  DFFQX1 \L12_reg[6]  ( .D(R11[6]), .CK(n59), .Q(L12[6]) );
  DFFQX1 \L12_reg[7]  ( .D(R11[7]), .CK(n55), .Q(L12[7]) );
  DFFQX1 \L12_reg[8]  ( .D(R11[8]), .CK(n14), .Q(L12[8]) );
  DFFQX1 \L12_reg[9]  ( .D(R11[9]), .CK(n3), .Q(L12[9]) );
  DFFQX1 \L12_reg[10]  ( .D(R11[10]), .CK(n76), .Q(L12[10]) );
  DFFQX1 \L12_reg[11]  ( .D(R11[11]), .CK(n75), .Q(L12[11]) );
  DFFQX1 \L12_reg[12]  ( .D(R11[12]), .CK(n74), .Q(L12[12]) );
  DFFQX1 \L12_reg[13]  ( .D(R11[13]), .CK(n73), .Q(L12[13]) );
  DFFQX1 \L12_reg[14]  ( .D(R11[14]), .CK(n69), .Q(L12[14]) );
  DFFQX1 \L12_reg[15]  ( .D(R11[15]), .CK(n68), .Q(L12[15]) );
  DFFQX1 \L12_reg[16]  ( .D(R11[16]), .CK(n88), .Q(L12[16]) );
  DFFQX1 \L12_reg[17]  ( .D(R11[17]), .CK(n18), .Q(L12[17]) );
  DFFQX1 \L12_reg[18]  ( .D(R11[18]), .CK(n17), .Q(L12[18]) );
  DFFQX1 \L12_reg[19]  ( .D(R11[19]), .CK(n16), .Q(L12[19]) );
  DFFQX1 \L12_reg[20]  ( .D(R11[20]), .CK(n12), .Q(L12[20]) );
  DFFQX1 \L12_reg[21]  ( .D(R11[21]), .CK(n11), .Q(L12[21]) );
  DFFQX1 \L12_reg[22]  ( .D(R11[22]), .CK(n10), .Q(L12[22]) );
  DFFQX1 \L12_reg[23]  ( .D(R11[23]), .CK(n9), .Q(L12[23]) );
  DFFQX1 \L12_reg[24]  ( .D(R11[24]), .CK(n5), .Q(L12[24]) );
  DFFQX1 \L12_reg[25]  ( .D(R11[25]), .CK(n4), .Q(L12[25]) );
  DFFQX1 \L12_reg[26]  ( .D(R11[26]), .CK(n25), .Q(L12[26]) );
  DFFQX1 \L12_reg[27]  ( .D(R11[27]), .CK(n24), .Q(L12[27]) );
  DFFQX1 \L12_reg[28]  ( .D(R11[28]), .CK(n23), .Q(L12[28]) );
  DFFQX1 \L12_reg[29]  ( .D(R11[29]), .CK(n102), .Q(L12[29]) );
  DFFQX1 \L12_reg[30]  ( .D(R11[30]), .CK(n99), .Q(L12[30]) );
  DFFQX1 \L12_reg[31]  ( .D(R11[31]), .CK(n101), .Q(L12[31]) );
  DFFQX1 \L12_reg[32]  ( .D(R11[32]), .CK(n119), .Q(L12[32]) );
  DFFQX1 \L13_reg[1]  ( .D(R12[1]), .CK(n136), .Q(L13[1]) );
  DFFQX1 \L13_reg[2]  ( .D(R12[2]), .CK(n128), .Q(L13[2]) );
  DFFQX1 \L13_reg[3]  ( .D(R12[3]), .CK(n142), .Q(L13[3]) );
  DFFQX1 \L13_reg[4]  ( .D(R12[4]), .CK(n119), .Q(L13[4]) );
  DFFQX1 \L13_reg[5]  ( .D(R12[5]), .CK(n101), .Q(L13[5]) );
  DFFQX1 \L13_reg[6]  ( .D(R12[6]), .CK(n104), .Q(L13[6]) );
  DFFQX1 \L13_reg[7]  ( .D(R12[7]), .CK(n133), .Q(L13[7]) );
  DFFQX1 \L13_reg[8]  ( .D(R12[8]), .CK(n140), .Q(L13[8]) );
  DFFQX1 \L13_reg[9]  ( .D(R12[9]), .CK(n132), .Q(L13[9]) );
  DFFQX1 \L13_reg[10]  ( .D(R12[10]), .CK(n131), .Q(L13[10]) );
  DFFQX1 \L13_reg[11]  ( .D(R12[11]), .CK(n130), .Q(L13[11]) );
  DFFQX1 \L13_reg[12]  ( .D(R12[12]), .CK(n141), .Q(L13[12]) );
  DFFQX1 \L13_reg[13]  ( .D(R12[13]), .CK(n137), .Q(L13[13]) );
  DFFQX1 \L13_reg[14]  ( .D(R12[14]), .CK(n85), .Q(L13[14]) );
  DFFQX1 \L13_reg[15]  ( .D(R12[15]), .CK(n93), .Q(L13[15]) );
  DFFQX1 \L13_reg[16]  ( .D(R12[16]), .CK(n125), .Q(L13[16]) );
  DFFQX1 \L13_reg[17]  ( .D(R12[17]), .CK(n126), .Q(L13[17]) );
  DFFQX1 \L13_reg[18]  ( .D(R12[18]), .CK(n22), .Q(L13[18]) );
  DFFQX1 \L13_reg[19]  ( .D(R12[19]), .CK(n127), .Q(L13[19]) );
  DFFQX1 \L13_reg[20]  ( .D(R12[20]), .CK(n78), .Q(L13[20]) );
  DFFQX1 \L13_reg[21]  ( .D(R12[21]), .CK(n98), .Q(L13[21]) );
  DFFQX1 \L13_reg[22]  ( .D(R12[22]), .CK(n104), .Q(L13[22]) );
  DFFQX1 \L13_reg[23]  ( .D(R12[23]), .CK(n139), .Q(L13[23]) );
  DFFQX1 \L13_reg[24]  ( .D(R12[24]), .CK(n123), .Q(L13[24]) );
  DFFQX1 \L13_reg[25]  ( .D(R12[25]), .CK(n114), .Q(L13[25]) );
  DFFQX1 \L13_reg[26]  ( .D(R12[26]), .CK(n115), .Q(L13[26]) );
  DFFQX1 \L13_reg[27]  ( .D(R12[27]), .CK(n116), .Q(L13[27]) );
  DFFQX1 \L13_reg[28]  ( .D(R12[28]), .CK(n117), .Q(L13[28]) );
  DFFQX1 \L13_reg[29]  ( .D(R12[29]), .CK(n118), .Q(L13[29]) );
  DFFQX1 \L13_reg[30]  ( .D(R12[30]), .CK(n121), .Q(L13[30]) );
  DFFQX1 \L13_reg[31]  ( .D(R12[31]), .CK(n122), .Q(L13[31]) );
  DFFQX1 \L13_reg[32]  ( .D(R12[32]), .CK(n103), .Q(L13[32]) );
  DFFQX1 \L14_reg[1]  ( .D(R13[1]), .CK(n125), .Q(L14[1]) );
  DFFQX1 \L14_reg[2]  ( .D(R13[2]), .CK(n126), .Q(L14[2]) );
  DFFQX1 \L14_reg[3]  ( .D(R13[3]), .CK(n57), .Q(L14[3]) );
  DFFQX1 \L14_reg[4]  ( .D(R13[4]), .CK(n127), .Q(L14[4]) );
  DFFQX1 \L14_reg[5]  ( .D(R13[5]), .CK(n98), .Q(L14[5]) );
  DFFQX1 \L14_reg[6]  ( .D(R13[6]), .CK(n138), .Q(L14[6]) );
  DFFQX1 \L14_reg[7]  ( .D(R13[7]), .CK(n144), .Q(L14[7]) );
  DFFQX1 \L14_reg[8]  ( .D(R13[8]), .CK(n97), .Q(L14[8]) );
  DFFQX1 \L14_reg[9]  ( .D(R13[9]), .CK(n101), .Q(L14[9]) );
  DFFQX1 \L14_reg[10]  ( .D(R13[10]), .CK(n119), .Q(L14[10]) );
  DFFQX1 \L14_reg[11]  ( .D(R13[11]), .CK(n99), .Q(L14[11]) );
  DFFQX1 \L14_reg[12]  ( .D(R13[12]), .CK(n100), .Q(L14[12]) );
  DFFQX1 \L14_reg[13]  ( .D(R13[13]), .CK(n102), .Q(L14[13]) );
  DFFQX1 \L14_reg[14]  ( .D(R13[14]), .CK(n143), .Q(L14[14]) );
  DFFQX1 \L14_reg[15]  ( .D(R13[15]), .CK(n132), .Q(L14[15]) );
  DFFQX1 \L14_reg[16]  ( .D(R13[16]), .CK(n130), .Q(L14[16]) );
  DFFQX1 \L14_reg[17]  ( .D(R13[17]), .CK(n137), .Q(L14[17]) );
  DFFQX1 \L14_reg[18]  ( .D(R13[18]), .CK(n135), .Q(L14[18]) );
  DFFQX1 \L14_reg[19]  ( .D(R13[19]), .CK(n140), .Q(L14[19]) );
  DFFQX1 \L14_reg[20]  ( .D(R13[20]), .CK(n141), .Q(L14[20]) );
  DFFQX1 \L14_reg[21]  ( .D(R13[21]), .CK(n121), .Q(L14[21]) );
  DFFQX1 \L14_reg[22]  ( .D(R13[22]), .CK(n142), .Q(L14[22]) );
  DFFQX1 \L14_reg[23]  ( .D(R13[23]), .CK(n27), .Q(L14[23]) );
  DFFQX1 \L14_reg[24]  ( .D(R13[24]), .CK(n129), .Q(L14[24]) );
  DFFQX1 \L14_reg[25]  ( .D(R13[25]), .CK(n131), .Q(L14[25]) );
  DFFQX1 \L14_reg[26]  ( .D(R13[26]), .CK(clk), .Q(L14[26]) );
  DFFQX1 \L14_reg[27]  ( .D(R13[27]), .CK(n136), .Q(L14[27]) );
  DFFQX1 \L14_reg[28]  ( .D(R13[28]), .CK(n94), .Q(L14[28]) );
  DFFQX1 \L14_reg[29]  ( .D(R13[29]), .CK(n134), .Q(L14[29]) );
  DFFQX1 \L14_reg[30]  ( .D(R13[30]), .CK(n133), .Q(L14[30]) );
  DFFQX1 \L14_reg[31]  ( .D(R13[31]), .CK(n139), .Q(L14[31]) );
  DFFQX1 \L14_reg[32]  ( .D(R13[32]), .CK(n128), .Q(L14[32]) );
  DFFQX1 \key_r_reg[50]  ( .D(key[50]), .CK(n96), .Q(key_r[50]) );
  DFFQX1 \key_r_reg[49]  ( .D(key[49]), .CK(n96), .Q(key_r[49]) );
  DFFQX1 \key_r_reg[46]  ( .D(key[46]), .CK(n96), .Q(key_r[46]) );
  DFFQX1 \key_r_reg[45]  ( .D(key[45]), .CK(n96), .Q(key_r[45]) );
  DFFQX1 \key_r_reg[43]  ( .D(key[43]), .CK(n96), .Q(key_r[43]) );
  DFFQX1 \key_r_reg[42]  ( .D(key[42]), .CK(n95), .Q(key_r[42]) );
  DFFQX1 \key_r_reg[39]  ( .D(key[39]), .CK(n95), .Q(key_r[39]) );
  DFFQX1 \key_r_reg[38]  ( .D(key[38]), .CK(n95), .Q(key_r[38]) );
  DFFQX1 \key_r_reg[18]  ( .D(key[18]), .CK(n93), .Q(key_r[18]) );
  DFFQX1 \key_r_reg[15]  ( .D(key[15]), .CK(n92), .Q(key_r[15]) );
  DFFQX1 \key_r_reg[12]  ( .D(key[12]), .CK(n92), .Q(key_r[12]) );
  DFFQX1 \key_r_reg[11]  ( .D(key[11]), .CK(n92), .Q(key_r[11]) );
  DFFQX1 \key_r_reg[10]  ( .D(key[10]), .CK(n92), .Q(key_r[10]) );
  DFFQX1 \key_r_reg[8]  ( .D(key[8]), .CK(n92), .Q(key_r[8]) );
  DFFQX1 \key_r_reg[5]  ( .D(key[5]), .CK(n91), .Q(key_r[5]) );
  DFFQX1 \key_r_reg[3]  ( .D(key[3]), .CK(n91), .Q(key_r[3]) );
  DFFQX1 \desIn_r_reg[55]  ( .D(desIn[55]), .CK(n90), .Q(desIn_r[55]) );
  DFFQX1 \desIn_r_reg[53]  ( .D(desIn[53]), .CK(n90), .Q(desIn_r[53]) );
  DFFQX1 \desIn_r_reg[51]  ( .D(desIn[51]), .CK(n89), .Q(desIn_r[51]) );
  DFFQX1 \desIn_r_reg[49]  ( .D(desIn[49]), .CK(n89), .Q(desIn_r[49]) );
  DFFQX1 \desIn_r_reg[47]  ( .D(desIn[47]), .CK(n89), .Q(desIn_r[47]) );
  DFFQX1 \desIn_r_reg[45]  ( .D(desIn[45]), .CK(n89), .Q(desIn_r[45]) );
  DFFQX1 \desIn_r_reg[43]  ( .D(desIn[43]), .CK(n88), .Q(desIn_r[43]) );
  DFFQX1 \desIn_r_reg[41]  ( .D(desIn[41]), .CK(n88), .Q(desIn_r[41]) );
  DFFQX1 \desIn_r_reg[23]  ( .D(desIn[23]), .CK(n86), .Q(desIn_r[23]) );
  DFFQX1 \desIn_r_reg[21]  ( .D(desIn[21]), .CK(n86), .Q(desIn_r[21]) );
  DFFQX1 \desIn_r_reg[19]  ( .D(desIn[19]), .CK(n86), .Q(desIn_r[19]) );
  DFFQX1 \desIn_r_reg[17]  ( .D(desIn[17]), .CK(n86), .Q(desIn_r[17]) );
  DFFQX1 \desIn_r_reg[15]  ( .D(desIn[15]), .CK(n85), .Q(desIn_r[15]) );
  DFFQX1 \desIn_r_reg[13]  ( .D(desIn[13]), .CK(n85), .Q(desIn_r[13]) );
  DFFQX1 \desIn_r_reg[11]  ( .D(desIn[11]), .CK(n85), .Q(desIn_r[11]) );
  DFFQX1 \desIn_r_reg[9]  ( .D(desIn[9]), .CK(n85), .Q(desIn_r[9]) );
  DFFQX1 \R0_reg[2]  ( .D(N1), .CK(n80), .Q(R0[2]) );
  DFFQX1 \R0_reg[3]  ( .D(N2), .CK(n80), .Q(R0[3]) );
  DFFQX1 \R0_reg[6]  ( .D(N5), .CK(n79), .Q(R0[6]) );
  DFFQX1 \R0_reg[7]  ( .D(N6), .CK(n79), .Q(R0[7]) );
  DFFQX1 \R0_reg[10]  ( .D(N9), .CK(n79), .Q(R0[10]) );
  DFFQX1 \R0_reg[11]  ( .D(N10), .CK(n79), .Q(R0[11]) );
  DFFQX1 \R0_reg[14]  ( .D(N13), .CK(n79), .Q(R0[14]) );
  DFFQX1 \R0_reg[15]  ( .D(N14), .CK(n78), .Q(R0[15]) );
  DFFQX1 \R0_reg[18]  ( .D(N17), .CK(n78), .Q(R0[18]) );
  DFFQX1 \R0_reg[19]  ( .D(N18), .CK(n78), .Q(R0[19]) );
  DFFQX1 \R0_reg[22]  ( .D(N21), .CK(n78), .Q(R0[22]) );
  DFFQX1 \R0_reg[23]  ( .D(N22), .CK(n78), .Q(R0[23]) );
  DFFQX1 \R0_reg[26]  ( .D(N25), .CK(n77), .Q(R0[26]) );
  DFFQX1 \R0_reg[27]  ( .D(N26), .CK(n77), .Q(R0[27]) );
  DFFQX1 \R0_reg[30]  ( .D(N29), .CK(n77), .Q(R0[30]) );
  DFFQX1 \R0_reg[31]  ( .D(N30), .CK(n77), .Q(R0[31]) );
  DFFQX1 \R1_reg[2]  ( .D(N33), .CK(n73), .Q(R1[2]) );
  DFFQX1 \R1_reg[3]  ( .D(N34), .CK(n73), .Q(R1[3]) );
  DFFQX1 \R1_reg[6]  ( .D(N37), .CK(n72), .Q(R1[6]) );
  DFFQX1 \R1_reg[7]  ( .D(N38), .CK(n72), .Q(R1[7]) );
  DFFQX1 \R1_reg[10]  ( .D(N41), .CK(n72), .Q(R1[10]) );
  DFFQX1 \R1_reg[11]  ( .D(N42), .CK(n72), .Q(R1[11]) );
  DFFQX1 \R1_reg[14]  ( .D(N45), .CK(n71), .Q(R1[14]) );
  DFFQX1 \R1_reg[15]  ( .D(N46), .CK(n71), .Q(R1[15]) );
  DFFQX1 \R1_reg[18]  ( .D(N49), .CK(n71), .Q(R1[18]) );
  DFFQX1 \R1_reg[19]  ( .D(N50), .CK(n71), .Q(R1[19]) );
  DFFQX1 \R1_reg[22]  ( .D(N53), .CK(n71), .Q(R1[22]) );
  DFFQX1 \R1_reg[23]  ( .D(N54), .CK(n70), .Q(R1[23]) );
  DFFQX1 \R1_reg[26]  ( .D(N57), .CK(n70), .Q(R1[26]) );
  DFFQX1 \R1_reg[27]  ( .D(N58), .CK(n70), .Q(R1[27]) );
  DFFQX1 \R1_reg[30]  ( .D(N61), .CK(n70), .Q(R1[30]) );
  DFFQX1 \R1_reg[31]  ( .D(N62), .CK(n70), .Q(R1[31]) );
  DFFQX1 \R2_reg[2]  ( .D(N65), .CK(n66), .Q(R2[2]) );
  DFFQX1 \R2_reg[3]  ( .D(N66), .CK(n66), .Q(R2[3]) );
  DFFQX1 \R2_reg[6]  ( .D(N69), .CK(n65), .Q(R2[6]) );
  DFFQX1 \R2_reg[7]  ( .D(N70), .CK(n65), .Q(R2[7]) );
  DFFQX1 \R2_reg[10]  ( .D(N73), .CK(n65), .Q(R2[10]) );
  DFFQX1 \R2_reg[11]  ( .D(N74), .CK(n65), .Q(R2[11]) );
  DFFQX1 \R2_reg[14]  ( .D(N77), .CK(n64), .Q(R2[14]) );
  DFFQX1 \R2_reg[15]  ( .D(N78), .CK(n64), .Q(R2[15]) );
  DFFQX1 \R2_reg[18]  ( .D(N81), .CK(n64), .Q(R2[18]) );
  DFFQX1 \R2_reg[19]  ( .D(N82), .CK(n64), .Q(R2[19]) );
  DFFQX1 \R2_reg[22]  ( .D(N85), .CK(n63), .Q(R2[22]) );
  DFFQX1 \R2_reg[23]  ( .D(N86), .CK(n63), .Q(R2[23]) );
  DFFQX1 \R2_reg[26]  ( .D(N89), .CK(n63), .Q(R2[26]) );
  DFFQX1 \R2_reg[27]  ( .D(N90), .CK(n63), .Q(R2[27]) );
  DFFQX1 \R2_reg[30]  ( .D(N93), .CK(n63), .Q(R2[30]) );
  DFFQX1 \R2_reg[31]  ( .D(N94), .CK(n62), .Q(R2[31]) );
  DFFQX1 \R3_reg[2]  ( .D(N97), .CK(n59), .Q(R3[2]) );
  DFFQX1 \R3_reg[3]  ( .D(N98), .CK(n58), .Q(R3[3]) );
  DFFQX1 \R3_reg[6]  ( .D(N101), .CK(n58), .Q(R3[6]) );
  DFFQX1 \R3_reg[7]  ( .D(N102), .CK(n58), .Q(R3[7]) );
  DFFQX1 \R3_reg[10]  ( .D(N105), .CK(n58), .Q(R3[10]) );
  DFFQX1 \R3_reg[11]  ( .D(N106), .CK(n58), .Q(R3[11]) );
  DFFQX1 \R3_reg[14]  ( .D(N109), .CK(n57), .Q(R3[14]) );
  DFFQX1 \R3_reg[15]  ( .D(N110), .CK(n57), .Q(R3[15]) );
  DFFQX1 \R3_reg[18]  ( .D(N113), .CK(n57), .Q(R3[18]) );
  DFFQX1 \R3_reg[19]  ( .D(N114), .CK(n57), .Q(R3[19]) );
  DFFQX1 \R3_reg[22]  ( .D(N117), .CK(n56), .Q(R3[22]) );
  DFFQX1 \R3_reg[23]  ( .D(N118), .CK(n56), .Q(R3[23]) );
  DFFQX1 \R3_reg[26]  ( .D(N121), .CK(n56), .Q(R3[26]) );
  DFFQX1 \R3_reg[27]  ( .D(N122), .CK(n56), .Q(R3[27]) );
  DFFQX1 \R3_reg[30]  ( .D(N125), .CK(n55), .Q(R3[30]) );
  DFFQX1 \R3_reg[31]  ( .D(N126), .CK(n55), .Q(R3[31]) );
  DFFQX1 \R4_reg[2]  ( .D(N129), .CK(n51), .Q(R4[2]) );
  DFFQX1 \R4_reg[3]  ( .D(N130), .CK(n51), .Q(R4[3]) );
  DFFQX1 \R4_reg[6]  ( .D(N133), .CK(n51), .Q(R4[6]) );
  DFFQX1 \R4_reg[7]  ( .D(N134), .CK(n51), .Q(R4[7]) );
  DFFQX1 \R4_reg[10]  ( .D(N137), .CK(n51), .Q(R4[10]) );
  DFFQX1 \R4_reg[11]  ( .D(N138), .CK(n50), .Q(R4[11]) );
  DFFQX1 \R4_reg[14]  ( .D(N141), .CK(n50), .Q(R4[14]) );
  DFFQX1 \R4_reg[15]  ( .D(N142), .CK(n50), .Q(R4[15]) );
  DFFQX1 \R4_reg[18]  ( .D(N145), .CK(n50), .Q(R4[18]) );
  DFFQX1 \R4_reg[19]  ( .D(N146), .CK(n50), .Q(R4[19]) );
  DFFQX1 \R4_reg[22]  ( .D(N149), .CK(n49), .Q(R4[22]) );
  DFFQX1 \R4_reg[23]  ( .D(N150), .CK(n49), .Q(R4[23]) );
  DFFQX1 \R4_reg[26]  ( .D(N153), .CK(n49), .Q(R4[26]) );
  DFFQX1 \R4_reg[27]  ( .D(N154), .CK(n49), .Q(R4[27]) );
  DFFQX1 \R4_reg[30]  ( .D(N157), .CK(n48), .Q(R4[30]) );
  DFFQX1 \R4_reg[31]  ( .D(N158), .CK(n48), .Q(R4[31]) );
  DFFQX1 \R5_reg[2]  ( .D(N161), .CK(n44), .Q(R5[2]) );
  DFFQX1 \R5_reg[3]  ( .D(N162), .CK(n44), .Q(R5[3]) );
  DFFQX1 \R5_reg[6]  ( .D(N165), .CK(n44), .Q(R5[6]) );
  DFFQX1 \R5_reg[7]  ( .D(N166), .CK(n44), .Q(R5[7]) );
  DFFQX1 \R5_reg[10]  ( .D(N169), .CK(n43), .Q(R5[10]) );
  DFFQX1 \R5_reg[11]  ( .D(N170), .CK(n43), .Q(R5[11]) );
  DFFQX1 \R5_reg[14]  ( .D(N173), .CK(n43), .Q(R5[14]) );
  DFFQX1 \R5_reg[15]  ( .D(N174), .CK(n43), .Q(R5[15]) );
  DFFQX1 \R5_reg[18]  ( .D(N177), .CK(n43), .Q(R5[18]) );
  DFFQX1 \R5_reg[19]  ( .D(N178), .CK(n42), .Q(R5[19]) );
  DFFQX1 \R5_reg[22]  ( .D(N181), .CK(n42), .Q(R5[22]) );
  DFFQX1 \R5_reg[23]  ( .D(N182), .CK(n42), .Q(R5[23]) );
  DFFQX1 \R5_reg[26]  ( .D(N185), .CK(n42), .Q(R5[26]) );
  DFFQX1 \R5_reg[27]  ( .D(N186), .CK(n42), .Q(R5[27]) );
  DFFQX1 \R5_reg[30]  ( .D(N189), .CK(n41), .Q(R5[30]) );
  DFFQX1 \R5_reg[31]  ( .D(N190), .CK(n41), .Q(R5[31]) );
  DFFQX1 \R6_reg[2]  ( .D(N193), .CK(n37), .Q(R6[2]) );
  DFFQX1 \R6_reg[3]  ( .D(N194), .CK(n37), .Q(R6[3]) );
  DFFQX1 \R6_reg[6]  ( .D(N197), .CK(n37), .Q(R6[6]) );
  DFFQX1 \R6_reg[7]  ( .D(N198), .CK(n37), .Q(R6[7]) );
  DFFQX1 \R6_reg[10]  ( .D(N201), .CK(n36), .Q(R6[10]) );
  DFFQX1 \R6_reg[11]  ( .D(N202), .CK(n36), .Q(R6[11]) );
  DFFQX1 \R6_reg[14]  ( .D(N205), .CK(n36), .Q(R6[14]) );
  DFFQX1 \R6_reg[15]  ( .D(N206), .CK(n36), .Q(R6[15]) );
  DFFQX1 \R6_reg[18]  ( .D(N209), .CK(n35), .Q(R6[18]) );
  DFFQX1 \R6_reg[19]  ( .D(N210), .CK(n35), .Q(R6[19]) );
  DFFQX1 \R6_reg[22]  ( .D(N213), .CK(n35), .Q(R6[22]) );
  DFFQX1 \R6_reg[23]  ( .D(N214), .CK(n35), .Q(R6[23]) );
  DFFQX1 \R6_reg[26]  ( .D(N217), .CK(n35), .Q(R6[26]) );
  DFFQX1 \R6_reg[27]  ( .D(N218), .CK(n34), .Q(R6[27]) );
  DFFQX1 \R6_reg[30]  ( .D(N221), .CK(n34), .Q(R6[30]) );
  DFFQX1 \R6_reg[31]  ( .D(N222), .CK(n34), .Q(R6[31]) );
  DFFQX1 \R7_reg[2]  ( .D(N225), .CK(n30), .Q(R7[2]) );
  DFFQX1 \R7_reg[3]  ( .D(N226), .CK(n30), .Q(R7[3]) );
  DFFQX1 \R7_reg[6]  ( .D(N229), .CK(n30), .Q(R7[6]) );
  DFFQX1 \R7_reg[7]  ( .D(N230), .CK(n30), .Q(R7[7]) );
  DFFQX1 \R7_reg[10]  ( .D(N233), .CK(n29), .Q(R7[10]) );
  DFFQX1 \R7_reg[11]  ( .D(N234), .CK(n29), .Q(R7[11]) );
  DFFQX1 \R7_reg[14]  ( .D(N237), .CK(n29), .Q(R7[14]) );
  DFFQX1 \R7_reg[15]  ( .D(N238), .CK(n29), .Q(R7[15]) );
  DFFQX1 \R7_reg[18]  ( .D(N241), .CK(n28), .Q(R7[18]) );
  DFFQX1 \R7_reg[19]  ( .D(N242), .CK(n28), .Q(R7[19]) );
  DFFQX1 \R7_reg[22]  ( .D(N245), .CK(n28), .Q(R7[22]) );
  DFFQX1 \R7_reg[23]  ( .D(N246), .CK(n28), .Q(R7[23]) );
  DFFQX1 \R7_reg[26]  ( .D(N249), .CK(n27), .Q(R7[26]) );
  DFFQX1 \R7_reg[27]  ( .D(N250), .CK(n27), .Q(R7[27]) );
  DFFQX1 \R7_reg[30]  ( .D(N253), .CK(n27), .Q(R7[30]) );
  DFFQX1 \R7_reg[31]  ( .D(N254), .CK(n27), .Q(R7[31]) );
  DFFQX1 \R8_reg[2]  ( .D(N257), .CK(n23), .Q(R8[2]) );
  DFFQX1 \R8_reg[3]  ( .D(N258), .CK(n23), .Q(R8[3]) );
  DFFQX1 \R8_reg[6]  ( .D(N261), .CK(n23), .Q(R8[6]) );
  DFFQX1 \R8_reg[7]  ( .D(N262), .CK(n22), .Q(R8[7]) );
  DFFQX1 \R8_reg[10]  ( .D(N265), .CK(n22), .Q(R8[10]) );
  DFFQX1 \R8_reg[11]  ( .D(N266), .CK(n22), .Q(R8[11]) );
  DFFQX1 \R8_reg[14]  ( .D(N269), .CK(n22), .Q(R8[14]) );
  DFFQX1 \R8_reg[15]  ( .D(N270), .CK(n22), .Q(R8[15]) );
  DFFQX1 \R8_reg[18]  ( .D(N273), .CK(n21), .Q(R8[18]) );
  DFFQX1 \R8_reg[19]  ( .D(N274), .CK(n21), .Q(R8[19]) );
  DFFQX1 \R8_reg[22]  ( .D(N277), .CK(n21), .Q(R8[22]) );
  DFFQX1 \R8_reg[23]  ( .D(N278), .CK(n21), .Q(R8[23]) );
  DFFQX1 \R8_reg[26]  ( .D(N281), .CK(n20), .Q(R8[26]) );
  DFFQX1 \R8_reg[27]  ( .D(N282), .CK(n20), .Q(R8[27]) );
  DFFQX1 \R8_reg[30]  ( .D(N285), .CK(n20), .Q(R8[30]) );
  DFFQX1 \R8_reg[31]  ( .D(N286), .CK(n20), .Q(R8[31]) );
  DFFQX1 \R9_reg[2]  ( .D(N289), .CK(n16), .Q(R9[2]) );
  DFFQX1 \R9_reg[3]  ( .D(N290), .CK(n16), .Q(R9[3]) );
  DFFQX1 \R9_reg[6]  ( .D(N293), .CK(n15), .Q(R9[6]) );
  DFFQX1 \R9_reg[7]  ( .D(N294), .CK(n15), .Q(R9[7]) );
  DFFQX1 \R9_reg[10]  ( .D(N297), .CK(n15), .Q(R9[10]) );
  DFFQX1 \R9_reg[11]  ( .D(N298), .CK(n15), .Q(R9[11]) );
  DFFQX1 \R9_reg[14]  ( .D(N301), .CK(n15), .Q(R9[14]) );
  DFFQX1 \R9_reg[15]  ( .D(N302), .CK(n14), .Q(R9[15]) );
  DFFQX1 \R9_reg[18]  ( .D(N305), .CK(n14), .Q(R9[18]) );
  DFFQX1 \R9_reg[19]  ( .D(N306), .CK(n14), .Q(R9[19]) );
  DFFQX1 \R9_reg[22]  ( .D(N309), .CK(n14), .Q(R9[22]) );
  DFFQX1 \R9_reg[23]  ( .D(N310), .CK(n14), .Q(R9[23]) );
  DFFQX1 \R9_reg[26]  ( .D(N313), .CK(n13), .Q(R9[26]) );
  DFFQX1 \R9_reg[27]  ( .D(N314), .CK(n13), .Q(R9[27]) );
  DFFQX1 \R9_reg[30]  ( .D(N317), .CK(n13), .Q(R9[30]) );
  DFFQX1 \R9_reg[31]  ( .D(N318), .CK(n13), .Q(R9[31]) );
  DFFQX1 \R10_reg[2]  ( .D(N321), .CK(n9), .Q(R10[2]) );
  DFFQX1 \R10_reg[3]  ( .D(N322), .CK(n9), .Q(R10[3]) );
  DFFQX1 \R10_reg[6]  ( .D(N325), .CK(n8), .Q(R10[6]) );
  DFFQX1 \R10_reg[7]  ( .D(N326), .CK(n8), .Q(R10[7]) );
  DFFQX1 \R10_reg[10]  ( .D(N329), .CK(n8), .Q(R10[10]) );
  DFFQX1 \R10_reg[11]  ( .D(N330), .CK(n8), .Q(R10[11]) );
  DFFQX1 \R10_reg[14]  ( .D(N333), .CK(n7), .Q(R10[14]) );
  DFFQX1 \R10_reg[15]  ( .D(N334), .CK(n7), .Q(R10[15]) );
  DFFQX1 \R10_reg[18]  ( .D(N337), .CK(n7), .Q(R10[18]) );
  DFFQX1 \R10_reg[19]  ( .D(N338), .CK(n7), .Q(R10[19]) );
  DFFQX1 \R10_reg[22]  ( .D(N341), .CK(n7), .Q(R10[22]) );
  DFFQX1 \R10_reg[23]  ( .D(N342), .CK(n6), .Q(R10[23]) );
  DFFQX1 \R10_reg[26]  ( .D(N345), .CK(n6), .Q(R10[26]) );
  DFFQX1 \R10_reg[27]  ( .D(N346), .CK(n6), .Q(R10[27]) );
  DFFQX1 \R10_reg[30]  ( .D(N349), .CK(n6), .Q(R10[30]) );
  DFFQX1 \R10_reg[31]  ( .D(N350), .CK(n6), .Q(R10[31]) );
  DFFQX1 \R11_reg[2]  ( .D(N353), .CK(n36), .Q(R11[2]) );
  DFFQX1 \R11_reg[3]  ( .D(N354), .CK(n2), .Q(R11[3]) );
  DFFQX1 \R11_reg[6]  ( .D(N357), .CK(n3), .Q(R11[6]) );
  DFFQX1 \R11_reg[7]  ( .D(N358), .CK(n3), .Q(R11[7]) );
  DFFQX1 \R11_reg[10]  ( .D(N361), .CK(n3), .Q(R11[10]) );
  DFFQX1 \R11_reg[11]  ( .D(N362), .CK(n3), .Q(R11[11]) );
  DFFQX1 \R11_reg[14]  ( .D(N365), .CK(n2), .Q(R11[14]) );
  DFFQX1 \R11_reg[15]  ( .D(N366), .CK(n2), .Q(R11[15]) );
  DFFQX1 \R11_reg[18]  ( .D(N369), .CK(n2), .Q(R11[18]) );
  DFFQX1 \R11_reg[19]  ( .D(N370), .CK(n2), .Q(R11[19]) );
  DFFQX1 \R11_reg[22]  ( .D(N373), .CK(n40), .Q(R11[22]) );
  DFFQX1 \R11_reg[23]  ( .D(N374), .CK(n39), .Q(R11[23]) );
  DFFQX1 \R11_reg[26]  ( .D(N377), .CK(n38), .Q(R11[26]) );
  DFFQX1 \R11_reg[27]  ( .D(N378), .CK(n33), .Q(R11[27]) );
  DFFQX1 \R11_reg[30]  ( .D(N381), .CK(n32), .Q(R11[30]) );
  DFFQX1 \R11_reg[31]  ( .D(N382), .CK(n54), .Q(R11[31]) );
  DFFQX1 \R12_reg[2]  ( .D(N385), .CK(n100), .Q(R12[2]) );
  DFFQX1 \R12_reg[3]  ( .D(N386), .CK(n51), .Q(R12[3]) );
  DFFQX1 \R12_reg[6]  ( .D(N389), .CK(n49), .Q(R12[6]) );
  DFFQX1 \R12_reg[7]  ( .D(N390), .CK(n48), .Q(R12[7]) );
  DFFQX1 \R12_reg[10]  ( .D(N393), .CK(n44), .Q(R12[10]) );
  DFFQX1 \R12_reg[11]  ( .D(N394), .CK(n42), .Q(R12[11]) );
  DFFQX1 \R12_reg[14]  ( .D(N397), .CK(n103), .Q(R12[14]) );
  DFFQX1 \R12_reg[15]  ( .D(N398), .CK(n125), .Q(R12[15]) );
  DFFQX1 \R12_reg[18]  ( .D(N401), .CK(n126), .Q(R12[18]) );
  DFFQX1 \R12_reg[19]  ( .D(N402), .CK(n29), .Q(R12[19]) );
  DFFQX1 \R12_reg[22]  ( .D(N405), .CK(n138), .Q(R12[22]) );
  DFFQX1 \R12_reg[23]  ( .D(N406), .CK(n144), .Q(R12[23]) );
  DFFQX1 \R12_reg[26]  ( .D(N409), .CK(n105), .Q(R12[26]) );
  DFFQX1 \R12_reg[27]  ( .D(N410), .CK(n106), .Q(R12[27]) );
  DFFQX1 \R12_reg[30]  ( .D(N413), .CK(n123), .Q(R12[30]) );
  DFFQX1 \R12_reg[31]  ( .D(N414), .CK(n124), .Q(R12[31]) );
  DFFQX1 \R13_reg[2]  ( .D(N417), .CK(n106), .Q(R13[2]) );
  DFFQX1 \R13_reg[3]  ( .D(N418), .CK(n107), .Q(R13[3]) );
  DFFQX1 \R13_reg[6]  ( .D(N421), .CK(n108), .Q(R13[6]) );
  DFFQX1 \R13_reg[7]  ( .D(N422), .CK(n109), .Q(R13[7]) );
  DFFQX1 \R13_reg[10]  ( .D(N425), .CK(n110), .Q(R13[10]) );
  DFFQX1 \R13_reg[11]  ( .D(N426), .CK(n113), .Q(R13[11]) );
  DFFQX1 \R13_reg[14]  ( .D(N429), .CK(n114), .Q(R13[14]) );
  DFFQX1 \R13_reg[15]  ( .D(N430), .CK(n115), .Q(R13[15]) );
  DFFQX1 \R13_reg[18]  ( .D(N433), .CK(n116), .Q(R13[18]) );
  DFFQX1 \R13_reg[19]  ( .D(N434), .CK(n117), .Q(R13[19]) );
  DFFQX1 \R13_reg[22]  ( .D(N437), .CK(n105), .Q(R13[22]) );
  DFFQX1 \R13_reg[23]  ( .D(N438), .CK(n106), .Q(R13[23]) );
  DFFQX1 \R13_reg[26]  ( .D(N441), .CK(n107), .Q(R13[26]) );
  DFFQX1 \R13_reg[27]  ( .D(N442), .CK(n108), .Q(R13[27]) );
  DFFQX1 \R13_reg[30]  ( .D(N445), .CK(n7), .Q(R13[30]) );
  DFFQX1 \R13_reg[31]  ( .D(N446), .CK(n52), .Q(R13[31]) );
  DFFQX1 \R14_reg[2]  ( .D(N449), .CK(n113), .Q(FP[34]) );
  DFFQX1 \R14_reg[3]  ( .D(N450), .CK(n114), .Q(FP[35]) );
  DFFQX1 \R14_reg[6]  ( .D(N453), .CK(n115), .Q(FP[38]) );
  DFFQX1 \R14_reg[7]  ( .D(N454), .CK(n116), .Q(FP[39]) );
  DFFQX1 \R14_reg[10]  ( .D(N457), .CK(n118), .Q(FP[42]) );
  DFFQX1 \R14_reg[11]  ( .D(N458), .CK(n142), .Q(FP[43]) );
  DFFQX1 \R14_reg[14]  ( .D(N461), .CK(n138), .Q(FP[46]) );
  DFFQX1 \R14_reg[15]  ( .D(N462), .CK(n143), .Q(FP[47]) );
  DFFQX1 \R14_reg[18]  ( .D(N465), .CK(n97), .Q(FP[50]) );
  DFFQX1 \R14_reg[19]  ( .D(N466), .CK(n135), .Q(FP[51]) );
  DFFQX1 \R14_reg[22]  ( .D(N469), .CK(n134), .Q(FP[54]) );
  DFFQX1 \R14_reg[23]  ( .D(N470), .CK(n133), .Q(FP[55]) );
  DFFQX1 \R14_reg[26]  ( .D(N473), .CK(n140), .Q(FP[58]) );
  DFFQX1 \R14_reg[27]  ( .D(N474), .CK(n132), .Q(FP[59]) );
  DFFQX1 \R14_reg[30]  ( .D(N477), .CK(n142), .Q(FP[62]) );
  DFFQX1 \R14_reg[31]  ( .D(N478), .CK(n144), .Q(FP[63]) );
  DFFQX1 \key_r_reg[4]  ( .D(key[4]), .CK(n91), .Q(key_r[4]) );
  DFFQX1 \key_r_reg[51]  ( .D(key[51]), .CK(n96), .Q(key_r[51]) );
  DFFQX1 \key_r_reg[48]  ( .D(key[48]), .CK(n96), .Q(key_r[48]) );
  DFFQX1 \key_r_reg[47]  ( .D(key[47]), .CK(n96), .Q(key_r[47]) );
  DFFQX1 \key_r_reg[44]  ( .D(key[44]), .CK(n96), .Q(key_r[44]) );
  DFFQX1 \key_r_reg[41]  ( .D(key[41]), .CK(n95), .Q(key_r[41]) );
  DFFQX1 \key_r_reg[37]  ( .D(key[37]), .CK(n95), .Q(key_r[37]) );
  DFFQX1 \key_r_reg[36]  ( .D(key[36]), .CK(n95), .Q(key_r[36]) );
  DFFQX1 \key_r_reg[35]  ( .D(key[35]), .CK(n95), .Q(key_r[35]) );
  DFFQX1 \key_r_reg[34]  ( .D(key[34]), .CK(n95), .Q(key_r[34]) );
  DFFQX1 \key_r_reg[33]  ( .D(key[33]), .CK(n94), .Q(key_r[33]) );
  DFFQX1 \key_r_reg[31]  ( .D(key[31]), .CK(n94), .Q(key_r[31]) );
  DFFQX1 \key_r_reg[28]  ( .D(key[28]), .CK(n94), .Q(key_r[28]) );
  DFFQX1 \key_r_reg[26]  ( .D(key[26]), .CK(n94), .Q(key_r[26]) );
  DFFQX1 \key_r_reg[25]  ( .D(key[25]), .CK(n94), .Q(key_r[25]) );
  DFFQX1 \key_r_reg[24]  ( .D(key[24]), .CK(n93), .Q(key_r[24]) );
  DFFQX1 \key_r_reg[23]  ( .D(key[23]), .CK(n93), .Q(key_r[23]) );
  DFFQX1 \key_r_reg[22]  ( .D(key[22]), .CK(n93), .Q(key_r[22]) );
  DFFQX1 \key_r_reg[21]  ( .D(key[21]), .CK(n93), .Q(key_r[21]) );
  DFFQX1 \key_r_reg[20]  ( .D(key[20]), .CK(n93), .Q(key_r[20]) );
  DFFQX1 \key_r_reg[19]  ( .D(key[19]), .CK(n93), .Q(key_r[19]) );
  DFFQX1 \key_r_reg[17]  ( .D(key[17]), .CK(n93), .Q(key_r[17]) );
  DFFQX1 \key_r_reg[16]  ( .D(key[16]), .CK(n93), .Q(key_r[16]) );
  DFFQX1 \key_r_reg[13]  ( .D(key[13]), .CK(n92), .Q(key_r[13]) );
  DFFQX1 \key_r_reg[9]  ( .D(key[9]), .CK(n92), .Q(key_r[9]) );
  DFFQX1 \key_r_reg[7]  ( .D(key[7]), .CK(n92), .Q(key_r[7]) );
  DFFQX1 \key_r_reg[6]  ( .D(key[6]), .CK(n91), .Q(key_r[6]) );
  DFFQX1 \key_r_reg[2]  ( .D(key[2]), .CK(n91), .Q(key_r[2]) );
  DFFQX1 \key_r_reg[0]  ( .D(key[0]), .CK(n91), .Q(key_r[0]) );
  DFFQX1 \key_r_reg[55]  ( .D(key[55]), .CK(n97), .Q(key_r[55]) );
  DFFQX1 \key_r_reg[54]  ( .D(key[54]), .CK(n97), .Q(key_r[54]) );
  DFFQX1 \key_r_reg[52]  ( .D(key[52]), .CK(n97), .Q(key_r[52]) );
  DFFQX1 \R0_reg[1]  ( .D(N0), .CK(n80), .Q(R0[1]) );
  DFFQX1 \R0_reg[4]  ( .D(N3), .CK(n80), .Q(R0[4]) );
  DFFQX1 \R0_reg[5]  ( .D(N4), .CK(n80), .Q(R0[5]) );
  DFFQX1 \R0_reg[9]  ( .D(N8), .CK(n79), .Q(R0[9]) );
  DFFQX1 \R0_reg[13]  ( .D(N12), .CK(n79), .Q(R0[13]) );
  DFFQX1 \R0_reg[17]  ( .D(N16), .CK(n78), .Q(R0[17]) );
  DFFQX1 \R0_reg[21]  ( .D(N20), .CK(n78), .Q(R0[21]) );
  DFFQX1 \R0_reg[24]  ( .D(N23), .CK(n77), .Q(R0[24]) );
  DFFQX1 \R0_reg[25]  ( .D(N24), .CK(n77), .Q(R0[25]) );
  DFFQX1 \R0_reg[28]  ( .D(N27), .CK(n77), .Q(R0[28]) );
  DFFQX1 \R0_reg[32]  ( .D(N31), .CK(n77), .Q(R0[32]) );
  DFFQX1 \R1_reg[1]  ( .D(N32), .CK(n73), .Q(R1[1]) );
  DFFQX1 \R1_reg[4]  ( .D(N35), .CK(n73), .Q(R1[4]) );
  DFFQX1 \R1_reg[5]  ( .D(N36), .CK(n72), .Q(R1[5]) );
  DFFQX1 \R1_reg[9]  ( .D(N40), .CK(n72), .Q(R1[9]) );
  DFFQX1 \R1_reg[13]  ( .D(N44), .CK(n72), .Q(R1[13]) );
  DFFQX1 \R1_reg[17]  ( .D(N48), .CK(n71), .Q(R1[17]) );
  DFFQX1 \R1_reg[21]  ( .D(N52), .CK(n71), .Q(R1[21]) );
  DFFQX1 \R1_reg[24]  ( .D(N55), .CK(n70), .Q(R1[24]) );
  DFFQX1 \R1_reg[25]  ( .D(N56), .CK(n70), .Q(R1[25]) );
  DFFQX1 \R1_reg[28]  ( .D(N59), .CK(n70), .Q(R1[28]) );
  DFFQX1 \R1_reg[32]  ( .D(N63), .CK(n69), .Q(R1[32]) );
  DFFQX1 \R2_reg[1]  ( .D(N64), .CK(n66), .Q(R2[1]) );
  DFFQX1 \R2_reg[4]  ( .D(N67), .CK(n65), .Q(R2[4]) );
  DFFQX1 \R2_reg[5]  ( .D(N68), .CK(n65), .Q(R2[5]) );
  DFFQX1 \R2_reg[9]  ( .D(N72), .CK(n65), .Q(R2[9]) );
  DFFQX1 \R2_reg[13]  ( .D(N76), .CK(n64), .Q(R2[13]) );
  DFFQX1 \R2_reg[17]  ( .D(N80), .CK(n64), .Q(R2[17]) );
  DFFQX1 \R2_reg[21]  ( .D(N84), .CK(n64), .Q(R2[21]) );
  DFFQX1 \R2_reg[24]  ( .D(N87), .CK(n63), .Q(R2[24]) );
  DFFQX1 \R2_reg[25]  ( .D(N88), .CK(n63), .Q(R2[25]) );
  DFFQX1 \R2_reg[28]  ( .D(N91), .CK(n63), .Q(R2[28]) );
  DFFQX1 \R2_reg[32]  ( .D(N95), .CK(n62), .Q(R2[32]) );
  DFFQX1 \R3_reg[1]  ( .D(N96), .CK(n59), .Q(R3[1]) );
  DFFQX1 \R3_reg[4]  ( .D(N99), .CK(n58), .Q(R3[4]) );
  DFFQX1 \R3_reg[5]  ( .D(N100), .CK(n58), .Q(R3[5]) );
  DFFQX1 \R3_reg[9]  ( .D(N104), .CK(n58), .Q(R3[9]) );
  DFFQX1 \R3_reg[13]  ( .D(N108), .CK(n57), .Q(R3[13]) );
  DFFQX1 \R3_reg[17]  ( .D(N112), .CK(n57), .Q(R3[17]) );
  DFFQX1 \R3_reg[21]  ( .D(N116), .CK(n56), .Q(R3[21]) );
  DFFQX1 \R3_reg[24]  ( .D(N119), .CK(n56), .Q(R3[24]) );
  DFFQX1 \R3_reg[25]  ( .D(N120), .CK(n56), .Q(R3[25]) );
  DFFQX1 \R3_reg[28]  ( .D(N123), .CK(n56), .Q(R3[28]) );
  DFFQX1 \R3_reg[32]  ( .D(N127), .CK(n55), .Q(R3[32]) );
  DFFQX1 \R4_reg[1]  ( .D(N128), .CK(n52), .Q(R4[1]) );
  DFFQX1 \R4_reg[4]  ( .D(N131), .CK(n51), .Q(R4[4]) );
  DFFQX1 \R4_reg[5]  ( .D(N132), .CK(n51), .Q(R4[5]) );
  DFFQX1 \R4_reg[9]  ( .D(N136), .CK(n51), .Q(R4[9]) );
  DFFQX1 \R4_reg[13]  ( .D(N140), .CK(n50), .Q(R4[13]) );
  DFFQX1 \R4_reg[17]  ( .D(N144), .CK(n50), .Q(R4[17]) );
  DFFQX1 \R4_reg[21]  ( .D(N148), .CK(n49), .Q(R4[21]) );
  DFFQX1 \R4_reg[24]  ( .D(N151), .CK(n49), .Q(R4[24]) );
  DFFQX1 \R4_reg[25]  ( .D(N152), .CK(n49), .Q(R4[25]) );
  DFFQX1 \R4_reg[28]  ( .D(N155), .CK(n49), .Q(R4[28]) );
  DFFQX1 \R4_reg[32]  ( .D(N159), .CK(n48), .Q(R4[32]) );
  DFFQX1 \R5_reg[1]  ( .D(N160), .CK(n44), .Q(R5[1]) );
  DFFQX1 \R5_reg[4]  ( .D(N163), .CK(n44), .Q(R5[4]) );
  DFFQX1 \R5_reg[5]  ( .D(N164), .CK(n44), .Q(R5[5]) );
  DFFQX1 \R5_reg[9]  ( .D(N168), .CK(n44), .Q(R5[9]) );
  DFFQX1 \R5_reg[13]  ( .D(N172), .CK(n43), .Q(R5[13]) );
  DFFQX1 \R5_reg[17]  ( .D(N176), .CK(n43), .Q(R5[17]) );
  DFFQX1 \R5_reg[21]  ( .D(N180), .CK(n42), .Q(R5[21]) );
  DFFQX1 \R5_reg[24]  ( .D(N183), .CK(n42), .Q(R5[24]) );
  DFFQX1 \R5_reg[25]  ( .D(N184), .CK(n42), .Q(R5[25]) );
  DFFQX1 \R5_reg[28]  ( .D(N187), .CK(n41), .Q(R5[28]) );
  DFFQX1 \R5_reg[32]  ( .D(N191), .CK(n41), .Q(R5[32]) );
  DFFQX1 \R6_reg[1]  ( .D(N192), .CK(n37), .Q(R6[1]) );
  DFFQX1 \R6_reg[4]  ( .D(N195), .CK(n37), .Q(R6[4]) );
  DFFQX1 \R6_reg[5]  ( .D(N196), .CK(n37), .Q(R6[5]) );
  DFFQX1 \R6_reg[9]  ( .D(N200), .CK(n36), .Q(R6[9]) );
  DFFQX1 \R6_reg[13]  ( .D(N204), .CK(n36), .Q(R6[13]) );
  DFFQX1 \R6_reg[17]  ( .D(N208), .CK(n36), .Q(R6[17]) );
  DFFQX1 \R6_reg[21]  ( .D(N212), .CK(n35), .Q(R6[21]) );
  DFFQX1 \R6_reg[24]  ( .D(N215), .CK(n35), .Q(R6[24]) );
  DFFQX1 \R6_reg[25]  ( .D(N216), .CK(n35), .Q(R6[25]) );
  DFFQX1 \R6_reg[28]  ( .D(N219), .CK(n34), .Q(R6[28]) );
  DFFQX1 \R6_reg[32]  ( .D(N223), .CK(n34), .Q(R6[32]) );
  DFFQX1 \R7_reg[1]  ( .D(N224), .CK(n30), .Q(R7[1]) );
  DFFQX1 \R7_reg[4]  ( .D(N227), .CK(n30), .Q(R7[4]) );
  DFFQX1 \R7_reg[5]  ( .D(N228), .CK(n30), .Q(R7[5]) );
  DFFQX1 \R7_reg[9]  ( .D(N232), .CK(n29), .Q(R7[9]) );
  DFFQX1 \R7_reg[13]  ( .D(N236), .CK(n29), .Q(R7[13]) );
  DFFQX1 \R7_reg[17]  ( .D(N240), .CK(n28), .Q(R7[17]) );
  DFFQX1 \R7_reg[21]  ( .D(N244), .CK(n28), .Q(R7[21]) );
  DFFQX1 \R7_reg[24]  ( .D(N247), .CK(n28), .Q(R7[24]) );
  DFFQX1 \R7_reg[25]  ( .D(N248), .CK(n28), .Q(R7[25]) );
  DFFQX1 \R7_reg[28]  ( .D(N251), .CK(n27), .Q(R7[28]) );
  DFFQX1 \R7_reg[32]  ( .D(N255), .CK(n27), .Q(R7[32]) );
  DFFQX1 \R8_reg[1]  ( .D(N256), .CK(n23), .Q(R8[1]) );
  DFFQX1 \R8_reg[4]  ( .D(N259), .CK(n23), .Q(R8[4]) );
  DFFQX1 \R8_reg[5]  ( .D(N260), .CK(n23), .Q(R8[5]) );
  DFFQX1 \R8_reg[9]  ( .D(N264), .CK(n22), .Q(R8[9]) );
  DFFQX1 \R8_reg[13]  ( .D(N268), .CK(n22), .Q(R8[13]) );
  DFFQX1 \R8_reg[17]  ( .D(N272), .CK(n21), .Q(R8[17]) );
  DFFQX1 \R8_reg[21]  ( .D(N276), .CK(n21), .Q(R8[21]) );
  DFFQX1 \R8_reg[24]  ( .D(N279), .CK(n21), .Q(R8[24]) );
  DFFQX1 \R8_reg[25]  ( .D(N280), .CK(n20), .Q(R8[25]) );
  DFFQX1 \R8_reg[28]  ( .D(N283), .CK(n20), .Q(R8[28]) );
  DFFQX1 \R8_reg[32]  ( .D(N287), .CK(n20), .Q(R8[32]) );
  DFFQX1 \R9_reg[1]  ( .D(N288), .CK(n16), .Q(R9[1]) );
  DFFQX1 \R9_reg[4]  ( .D(N291), .CK(n16), .Q(R9[4]) );
  DFFQX1 \R9_reg[5]  ( .D(N292), .CK(n16), .Q(R9[5]) );
  DFFQX1 \R9_reg[9]  ( .D(N296), .CK(n15), .Q(R9[9]) );
  DFFQX1 \R9_reg[13]  ( .D(N300), .CK(n15), .Q(R9[13]) );
  DFFQX1 \R9_reg[17]  ( .D(N304), .CK(n14), .Q(R9[17]) );
  DFFQX1 \R9_reg[21]  ( .D(N308), .CK(n14), .Q(R9[21]) );
  DFFQX1 \R9_reg[24]  ( .D(N311), .CK(n13), .Q(R9[24]) );
  DFFQX1 \R9_reg[25]  ( .D(N312), .CK(n13), .Q(R9[25]) );
  DFFQX1 \R9_reg[28]  ( .D(N315), .CK(n13), .Q(R9[28]) );
  DFFQX1 \R9_reg[32]  ( .D(N319), .CK(n13), .Q(R9[32]) );
  DFFQX1 \R10_reg[1]  ( .D(N320), .CK(n9), .Q(R10[1]) );
  DFFQX1 \R10_reg[4]  ( .D(N323), .CK(n9), .Q(R10[4]) );
  DFFQX1 \R10_reg[5]  ( .D(N324), .CK(n8), .Q(R10[5]) );
  DFFQX1 \R10_reg[9]  ( .D(N328), .CK(n8), .Q(R10[9]) );
  DFFQX1 \R10_reg[13]  ( .D(N332), .CK(n8), .Q(R10[13]) );
  DFFQX1 \R10_reg[17]  ( .D(N336), .CK(n7), .Q(R10[17]) );
  DFFQX1 \R10_reg[21]  ( .D(N340), .CK(n7), .Q(R10[21]) );
  DFFQX1 \R10_reg[24]  ( .D(N343), .CK(n6), .Q(R10[24]) );
  DFFQX1 \R10_reg[25]  ( .D(N344), .CK(n6), .Q(R10[25]) );
  DFFQX1 \R10_reg[28]  ( .D(N347), .CK(n6), .Q(R10[28]) );
  DFFQX1 \R10_reg[32]  ( .D(N351), .CK(n5), .Q(R10[32]) );
  DFFQX1 \R11_reg[1]  ( .D(N352), .CK(n91), .Q(R11[1]) );
  DFFQX1 \R11_reg[4]  ( .D(N355), .CK(n3), .Q(R11[4]) );
  DFFQX1 \R11_reg[5]  ( .D(N356), .CK(n3), .Q(R11[5]) );
  DFFQX1 \R11_reg[9]  ( .D(N360), .CK(n3), .Q(R11[9]) );
  DFFQX1 \R11_reg[13]  ( .D(N364), .CK(n2), .Q(R11[13]) );
  DFFQX1 \R11_reg[17]  ( .D(N368), .CK(n2), .Q(R11[17]) );
  DFFQX1 \R11_reg[21]  ( .D(N372), .CK(n2), .Q(R11[21]) );
  DFFQX1 \R11_reg[24]  ( .D(N375), .CK(n31), .Q(R11[24]) );
  DFFQX1 \R11_reg[25]  ( .D(N376), .CK(n30), .Q(R11[25]) );
  DFFQX1 \R11_reg[28]  ( .D(N379), .CK(n26), .Q(R11[28]) );
  DFFQX1 \R11_reg[32]  ( .D(N383), .CK(n89), .Q(R11[32]) );
  DFFQX1 \R12_reg[1]  ( .D(N384), .CK(n100), .Q(R12[1]) );
  DFFQX1 \R12_reg[4]  ( .D(N387), .CK(n41), .Q(R12[4]) );
  DFFQX1 \R12_reg[5]  ( .D(N388), .CK(n37), .Q(R12[5]) );
  DFFQX1 \R12_reg[9]  ( .D(N392), .CK(n35), .Q(R12[9]) );
  DFFQX1 \R12_reg[13]  ( .D(N396), .CK(n127), .Q(R12[13]) );
  DFFQX1 \R12_reg[17]  ( .D(N400), .CK(n79), .Q(R12[17]) );
  DFFQX1 \R12_reg[21]  ( .D(N404), .CK(n107), .Q(R12[21]) );
  DFFQX1 \R12_reg[24]  ( .D(N407), .CK(n108), .Q(R12[24]) );
  DFFQX1 \R12_reg[25]  ( .D(N408), .CK(n109), .Q(R12[25]) );
  DFFQX1 \R12_reg[28]  ( .D(N411), .CK(n110), .Q(R12[28]) );
  DFFQX1 \R12_reg[32]  ( .D(N415), .CK(n129), .Q(R12[32]) );
  DFFQX1 \R13_reg[1]  ( .D(N416), .CK(n124), .Q(R13[1]) );
  DFFQX1 \R13_reg[4]  ( .D(N419), .CK(n111), .Q(R13[4]) );
  DFFQX1 \R13_reg[5]  ( .D(N420), .CK(n112), .Q(R13[5]) );
  DFFQX1 \R13_reg[9]  ( .D(N424), .CK(n113), .Q(R13[9]) );
  DFFQX1 \R13_reg[13]  ( .D(N428), .CK(n118), .Q(R13[13]) );
  DFFQX1 \R13_reg[17]  ( .D(N432), .CK(n121), .Q(R13[17]) );
  DFFQX1 \R13_reg[21]  ( .D(N436), .CK(n109), .Q(R13[21]) );
  DFFQX1 \R13_reg[24]  ( .D(N439), .CK(n110), .Q(R13[24]) );
  DFFQX1 \R13_reg[25]  ( .D(N440), .CK(n111), .Q(R13[25]) );
  DFFQX1 \R13_reg[28]  ( .D(N443), .CK(n112), .Q(R13[28]) );
  DFFQX1 \R13_reg[32]  ( .D(N447), .CK(n96), .Q(R13[32]) );
  DFFQX1 \R14_reg[1]  ( .D(N448), .CK(n122), .Q(FP[33]) );
  DFFQX1 \R14_reg[4]  ( .D(N451), .CK(n134), .Q(FP[36]) );
  DFFQX1 \R14_reg[5]  ( .D(N452), .CK(n105), .Q(FP[37]) );
  DFFQX1 \R14_reg[9]  ( .D(N456), .CK(n143), .Q(FP[41]) );
  DFFQX1 \R14_reg[13]  ( .D(N460), .CK(n99), .Q(FP[45]) );
  DFFQX1 \R14_reg[17]  ( .D(N464), .CK(n100), .Q(FP[49]) );
  DFFQX1 \R14_reg[21]  ( .D(N468), .CK(n131), .Q(FP[53]) );
  DFFQX1 \R14_reg[24]  ( .D(N471), .CK(n130), .Q(FP[56]) );
  DFFQX1 \R14_reg[25]  ( .D(N472), .CK(n141), .Q(FP[57]) );
  DFFQX1 \R14_reg[28]  ( .D(N475), .CK(n143), .Q(FP[60]) );
  DFFQX1 \R14_reg[32]  ( .D(N479), .CK(n102), .Q(FP[64]) );
  DFFQX1 \key_r_reg[40]  ( .D(key[40]), .CK(n95), .Q(key_r[40]) );
  DFFQX1 \key_r_reg[53]  ( .D(key[53]), .CK(n97), .Q(key_r[53]) );
  DFFQX1 \key_r_reg[32]  ( .D(key[32]), .CK(n94), .Q(key_r[32]) );
  DFFQX1 \key_r_reg[30]  ( .D(key[30]), .CK(n94), .Q(key_r[30]) );
  DFFQX1 \key_r_reg[29]  ( .D(key[29]), .CK(n94), .Q(key_r[29]) );
  DFFQX1 \key_r_reg[27]  ( .D(key[27]), .CK(n94), .Q(key_r[27]) );
  DFFQX1 \key_r_reg[14]  ( .D(key[14]), .CK(n92), .Q(key_r[14]) );
  DFFQX1 \key_r_reg[1]  ( .D(key[1]), .CK(n91), .Q(key_r[1]) );
  DFFQX1 \desIn_r_reg[59]  ( .D(desIn[59]), .CK(n90), .Q(desIn_r[59]) );
  DFFQX1 \desIn_r_reg[57]  ( .D(desIn[57]), .CK(n90), .Q(desIn_r[57]) );
  DFFQX1 \desIn_r_reg[39]  ( .D(desIn[39]), .CK(n88), .Q(desIn_r[39]) );
  DFFQX1 \desIn_r_reg[37]  ( .D(desIn[37]), .CK(n88), .Q(desIn_r[37]) );
  DFFQX1 \desIn_r_reg[35]  ( .D(desIn[35]), .CK(n88), .Q(desIn_r[35]) );
  DFFQX1 \desIn_r_reg[31]  ( .D(desIn[31]), .CK(n87), .Q(desIn_r[31]) );
  DFFQX1 \desIn_r_reg[25]  ( .D(desIn[25]), .CK(n86), .Q(desIn_r[25]) );
  DFFQX1 \desIn_r_reg[7]  ( .D(desIn[7]), .CK(n84), .Q(desIn_r[7]) );
  DFFQX1 \desIn_r_reg[5]  ( .D(desIn[5]), .CK(n84), .Q(desIn_r[5]) );
  DFFQX1 \desIn_r_reg[3]  ( .D(desIn[3]), .CK(n84), .Q(desIn_r[3]) );
  DFFQX1 \desIn_r_reg[1]  ( .D(desIn[1]), .CK(n84), .Q(desIn_r[1]) );
  DFFQX2 \R13_reg[20]  ( .D(N435), .CK(n124), .Q(R13[20]) );
  DFFQX2 \R10_reg[20]  ( .D(N339), .CK(n7), .Q(R10[20]) );
  DFFQX2 \R9_reg[20]  ( .D(N307), .CK(n14), .Q(R9[20]) );
  DFFQX2 \R8_reg[20]  ( .D(N275), .CK(n21), .Q(R8[20]) );
  DFFQX2 \R7_reg[20]  ( .D(N243), .CK(n28), .Q(R7[20]) );
  DFFQX2 \R6_reg[20]  ( .D(N211), .CK(n35), .Q(R6[20]) );
  DFFQX2 \R5_reg[20]  ( .D(N179), .CK(n42), .Q(R5[20]) );
  DFFQX2 \R4_reg[20]  ( .D(N147), .CK(n49), .Q(R4[20]) );
  DFFQX2 \R3_reg[20]  ( .D(N115), .CK(n57), .Q(R3[20]) );
  DFFQX2 \R2_reg[20]  ( .D(N83), .CK(n64), .Q(R2[20]) );
  DFFQX2 \desIn_r_reg[27]  ( .D(desIn[27]), .CK(n87), .Q(desIn_r[27]) );
  DFFQX2 \R7_reg[29]  ( .D(N252), .CK(n27), .Q(R7[29]) );
  DFFQX2 \R2_reg[29]  ( .D(N92), .CK(n63), .Q(R2[29]) );
  DFFQX2 \R11_reg[20]  ( .D(N371), .CK(n2), .Q(R11[20]) );
  DFFQX2 \R12_reg[12]  ( .D(N395), .CK(n45), .Q(R12[12]) );
  DFFQX2 \R14_reg[12]  ( .D(N459), .CK(n101), .Q(FP[44]) );
  DFFQX2 \R13_reg[12]  ( .D(N427), .CK(n104), .Q(R13[12]) );
  DFFQX2 \R11_reg[12]  ( .D(N363), .CK(n3), .Q(R11[12]) );
  DFFQX2 \R9_reg[12]  ( .D(N299), .CK(n15), .Q(R9[12]) );
  DFFQX2 \R8_reg[12]  ( .D(N267), .CK(n22), .Q(R8[12]) );
  DFFQX2 \R7_reg[12]  ( .D(N235), .CK(n29), .Q(R7[12]) );
  DFFQX2 \R5_reg[12]  ( .D(N171), .CK(n43), .Q(R5[12]) );
  DFFQX2 \R4_reg[12]  ( .D(N139), .CK(n50), .Q(R4[12]) );
  DFFQX2 \R3_reg[12]  ( .D(N107), .CK(n57), .Q(R3[12]) );
  DFFQX2 \R2_reg[12]  ( .D(N75), .CK(n65), .Q(R2[12]) );
  DFFQX2 \R0_reg[12]  ( .D(N11), .CK(n79), .Q(R0[12]) );
  DFFQX2 \desIn_r_reg[29]  ( .D(desIn[29]), .CK(n87), .Q(desIn_r[29]) );
  DFFQX2 \R6_reg[16]  ( .D(N207), .CK(n36), .Q(R6[16]) );
  DFFQX2 \R12_reg[20]  ( .D(N403), .CK(n19), .Q(R12[20]) );
  DFFQX2 \R1_reg[20]  ( .D(N51), .CK(n71), .Q(R1[20]) );
  DFFQX2 \R14_reg[20]  ( .D(N467), .CK(n139), .Q(FP[52]) );
  DFFQX2 \R0_reg[20]  ( .D(N19), .CK(n78), .Q(R0[20]) );
  DFFQX2 \R7_reg[8]  ( .D(N231), .CK(n29), .Q(R7[8]) );
  DFFQX2 \R2_reg[8]  ( .D(N71), .CK(n65), .Q(R2[8]) );
  DFFQX2 \R12_reg[29]  ( .D(N412), .CK(n97), .Q(R12[29]) );
  DFFQX2 \R1_reg[29]  ( .D(N60), .CK(n70), .Q(R1[29]) );
  DFFQX2 \R14_reg[29]  ( .D(N476), .CK(n119), .Q(FP[61]) );
  DFFQX2 \R13_reg[29]  ( .D(N444), .CK(n129), .Q(R13[29]) );
  DFFQX2 \R11_reg[29]  ( .D(N380), .CK(n46), .Q(R11[29]) );
  DFFQX2 \R10_reg[29]  ( .D(N348), .CK(n6), .Q(R10[29]) );
  DFFQX2 \R9_reg[29]  ( .D(N316), .CK(n13), .Q(R9[29]) );
  DFFQX2 \R6_reg[29]  ( .D(N220), .CK(n34), .Q(R6[29]) );
  DFFQX2 \R5_reg[29]  ( .D(N188), .CK(n41), .Q(R5[29]) );
  DFFQX2 \R4_reg[29]  ( .D(N156), .CK(n48), .Q(R4[29]) );
  DFFQX2 \R3_reg[29]  ( .D(N124), .CK(n56), .Q(R3[29]) );
  DFFQX2 \R0_reg[29]  ( .D(N28), .CK(n77), .Q(R0[29]) );
  DFFQX2 \desIn_r_reg[33]  ( .D(desIn[33]), .CK(n87), .Q(desIn_r[33]) );
  DFFQX2 \R12_reg[16]  ( .D(N399), .CK(n99), .Q(R12[16]) );
  DFFQX2 \R1_reg[16]  ( .D(N47), .CK(n71), .Q(R1[16]) );
  DFFQX2 \R14_reg[16]  ( .D(N463), .CK(n84), .Q(FP[48]) );
  DFFQX2 \R13_reg[16]  ( .D(N431), .CK(n123), .Q(R13[16]) );
  DFFQX2 \R11_reg[16]  ( .D(N367), .CK(n2), .Q(R11[16]) );
  DFFQX2 \R10_reg[16]  ( .D(N335), .CK(n7), .Q(R10[16]) );
  DFFQX2 \R9_reg[16]  ( .D(N303), .CK(n14), .Q(R9[16]) );
  DFFQX2 \R8_reg[16]  ( .D(N271), .CK(n21), .Q(R8[16]) );
  DFFQX2 \R7_reg[16]  ( .D(N239), .CK(n29), .Q(R7[16]) );
  DFFQX2 \R5_reg[16]  ( .D(N175), .CK(n43), .Q(R5[16]) );
  DFFQX2 \R4_reg[16]  ( .D(N143), .CK(n50), .Q(R4[16]) );
  DFFQX2 \R3_reg[16]  ( .D(N111), .CK(n57), .Q(R3[16]) );
  DFFQX2 \R2_reg[16]  ( .D(N79), .CK(n64), .Q(R2[16]) );
  DFFQX2 \R0_reg[16]  ( .D(N15), .CK(n78), .Q(R0[16]) );
  DFFQX2 \desIn_r_reg[61]  ( .D(desIn[61]), .CK(n90), .Q(desIn_r[61]) );
  DFFQX2 \R12_reg[8]  ( .D(N391), .CK(n34), .Q(R12[8]) );
  DFFQX2 \R14_reg[8]  ( .D(N455), .CK(n143), .Q(FP[40]) );
  DFFQX2 \R13_reg[8]  ( .D(N423), .CK(n142), .Q(R13[8]) );
  DFFQX2 \R11_reg[8]  ( .D(N359), .CK(n3), .Q(R11[8]) );
  DFFQX2 \R10_reg[8]  ( .D(N327), .CK(n8), .Q(R10[8]) );
  DFFQX2 \R9_reg[8]  ( .D(N295), .CK(n15), .Q(R9[8]) );
  DFFQX2 \R8_reg[8]  ( .D(N263), .CK(n22), .Q(R8[8]) );
  DFFQX2 \R6_reg[8]  ( .D(N199), .CK(n37), .Q(R6[8]) );
  DFFQX2 \R5_reg[8]  ( .D(N167), .CK(n44), .Q(R5[8]) );
  DFFQX2 \R4_reg[8]  ( .D(N135), .CK(n51), .Q(R4[8]) );
  DFFQX2 \R3_reg[8]  ( .D(N103), .CK(n58), .Q(R3[8]) );
  DFFQX2 \R0_reg[8]  ( .D(N7), .CK(n79), .Q(R0[8]) );
  DFFQX2 \R8_reg[29]  ( .D(N284), .CK(n20), .Q(R8[29]) );
  DFFQX2 \R1_reg[12]  ( .D(N43), .CK(n72), .Q(R1[12]) );
  DFFQX2 \R10_reg[12]  ( .D(N331), .CK(n8), .Q(R10[12]) );
  DFFQX2 \R6_reg[12]  ( .D(N203), .CK(n36), .Q(R6[12]) );
  DFFQX2 \R1_reg[8]  ( .D(N39), .CK(n72), .Q(R1[8]) );
  DFFQX2 \desIn_r_reg[63]  ( .D(desIn[63]), .CK(n91), .Q(desIn_r[63]) );
  CLKBUFX4 U3 ( .A(n111), .Y(n56) );
  CLKBUFX4 U4 ( .A(n111), .Y(n58) );
  CLKBUFX4 U5 ( .A(n109), .Y(n63) );
  CLKBUFX4 U6 ( .A(n107), .Y(n70) );
  CLKBUFX4 U7 ( .A(n138), .Y(n2) );
  CLKBUFX4 U8 ( .A(n118), .Y(n36) );
  CLKBUFX4 U9 ( .A(n116), .Y(n43) );
  CLKBUFX4 U10 ( .A(n113), .Y(n50) );
  CLKBUFX4 U11 ( .A(n104), .Y(n78) );
  CLKBUFX4 U12 ( .A(n104), .Y(n79) );
  CLKBUFX4 U13 ( .A(n127), .Y(n7) );
  CLKBUFX4 U14 ( .A(n21), .Y(n8) );
  CLKBUFX4 U15 ( .A(n120), .Y(n29) );
  CLKBUFX4 U16 ( .A(n111), .Y(n57) );
  CLKBUFX4 U17 ( .A(n125), .Y(n15) );
  CLKBUFX4 U18 ( .A(n122), .Y(n23) );
  CLKBUFX4 U19 ( .A(n122), .Y(n24) );
  CLKBUFX4 U20 ( .A(n122), .Y(n25) );
  CLKBUFX4 U21 ( .A(n121), .Y(n26) );
  CLKBUFX4 U22 ( .A(n120), .Y(n30) );
  CLKBUFX4 U23 ( .A(n120), .Y(n31) );
  CLKBUFX4 U24 ( .A(n119), .Y(n32) );
  CLKBUFX4 U25 ( .A(n115), .Y(n45) );
  CLKBUFX4 U26 ( .A(n115), .Y(n46) );
  CLKBUFX4 U27 ( .A(n114), .Y(n47) );
  CLKBUFX4 U28 ( .A(n113), .Y(n52) );
  CLKBUFX4 U29 ( .A(n112), .Y(n54) );
  CLKBUFX4 U30 ( .A(n112), .Y(n55) );
  CLKBUFX4 U31 ( .A(n110), .Y(n59) );
  CLKBUFX4 U32 ( .A(n110), .Y(n60) );
  CLKBUFX4 U33 ( .A(n107), .Y(n68) );
  CLKBUFX4 U34 ( .A(n107), .Y(n69) );
  CLKBUFX4 U35 ( .A(n106), .Y(n73) );
  CLKBUFX4 U36 ( .A(n105), .Y(n74) );
  CLKBUFX4 U37 ( .A(n92), .Y(n4) );
  CLKBUFX4 U38 ( .A(n127), .Y(n5) );
  CLKBUFX4 U39 ( .A(n15), .Y(n9) );
  CLKBUFX4 U40 ( .A(n124), .Y(n19) );
  CLKBUFX4 U41 ( .A(n98), .Y(n95) );
  CLKBUFX4 U42 ( .A(n98), .Y(n96) );
  CLKBUFX4 U43 ( .A(n99), .Y(n92) );
  CLKBUFX4 U44 ( .A(n99), .Y(n93) );
  CLKBUFX4 U45 ( .A(n121), .Y(n27) );
  CLKBUFX4 U46 ( .A(n121), .Y(n28) );
  CLKBUFX4 U47 ( .A(n103), .Y(n82) );
  CLKBUFX4 U48 ( .A(n119), .Y(n34) );
  CLKBUFX4 U49 ( .A(n118), .Y(n35) );
  CLKBUFX4 U50 ( .A(n118), .Y(n37) );
  BUFX4 U51 ( .A(n102), .Y(n3) );
  BUFX4 U52 ( .A(n127), .Y(n6) );
  BUFX4 U53 ( .A(n128), .Y(n10) );
  BUFX4 U54 ( .A(n126), .Y(n11) );
  BUFX4 U55 ( .A(n126), .Y(n12) );
  BUFX4 U56 ( .A(n126), .Y(n13) );
  BUFX4 U57 ( .A(n125), .Y(n14) );
  BUFX4 U58 ( .A(n125), .Y(n16) );
  BUFX4 U59 ( .A(n124), .Y(n17) );
  BUFX4 U60 ( .A(n124), .Y(n18) );
  BUFX4 U61 ( .A(n123), .Y(n20) );
  BUFX4 U62 ( .A(n123), .Y(n21) );
  BUFX4 U63 ( .A(n123), .Y(n22) );
  BUFX4 U64 ( .A(n119), .Y(n33) );
  BUFX4 U65 ( .A(n117), .Y(n38) );
  BUFX4 U66 ( .A(n117), .Y(n39) );
  BUFX4 U67 ( .A(n117), .Y(n40) );
  BUFX4 U68 ( .A(n116), .Y(n41) );
  BUFX4 U69 ( .A(n116), .Y(n42) );
  BUFX4 U70 ( .A(n115), .Y(n44) );
  BUFX4 U71 ( .A(n114), .Y(n48) );
  BUFX4 U72 ( .A(n114), .Y(n49) );
  BUFX4 U73 ( .A(n113), .Y(n51) );
  BUFX4 U74 ( .A(n112), .Y(n53) );
  BUFX4 U75 ( .A(n110), .Y(n61) );
  BUFX4 U76 ( .A(n109), .Y(n62) );
  BUFX4 U77 ( .A(n109), .Y(n64) );
  BUFX4 U78 ( .A(n108), .Y(n65) );
  BUFX4 U79 ( .A(n108), .Y(n66) );
  BUFX4 U80 ( .A(n108), .Y(n67) );
  BUFX4 U81 ( .A(n106), .Y(n71) );
  BUFX4 U82 ( .A(n106), .Y(n72) );
  BUFX4 U83 ( .A(n105), .Y(n75) );
  BUFX4 U84 ( .A(n105), .Y(n76) );
  BUFX4 U85 ( .A(n104), .Y(n77) );
  BUFX4 U86 ( .A(n103), .Y(n80) );
  BUFX4 U87 ( .A(n103), .Y(n81) );
  BUFX4 U88 ( .A(n102), .Y(n83) );
  BUFX4 U89 ( .A(n102), .Y(n84) );
  BUFX4 U90 ( .A(n102), .Y(n85) );
  BUFX4 U91 ( .A(n101), .Y(n86) );
  BUFX4 U92 ( .A(n101), .Y(n87) );
  BUFX4 U93 ( .A(n101), .Y(n88) );
  BUFX4 U94 ( .A(n100), .Y(n89) );
  BUFX4 U95 ( .A(n100), .Y(n90) );
  BUFX4 U96 ( .A(n100), .Y(n91) );
  BUFX4 U97 ( .A(n99), .Y(n94) );
  CLKBUFX3 U98 ( .A(n128), .Y(n127) );
  CLKBUFX3 U99 ( .A(n128), .Y(n126) );
  CLKBUFX3 U100 ( .A(n129), .Y(n125) );
  CLKBUFX3 U101 ( .A(n129), .Y(n124) );
  CLKBUFX3 U102 ( .A(n129), .Y(n123) );
  CLKBUFX3 U103 ( .A(n130), .Y(n122) );
  CLKBUFX3 U104 ( .A(n130), .Y(n121) );
  CLKBUFX3 U105 ( .A(n130), .Y(n120) );
  CLKBUFX3 U106 ( .A(n131), .Y(n119) );
  CLKBUFX3 U107 ( .A(n131), .Y(n118) );
  CLKBUFX3 U108 ( .A(n131), .Y(n117) );
  CLKBUFX3 U109 ( .A(n132), .Y(n116) );
  CLKBUFX3 U110 ( .A(n132), .Y(n115) );
  CLKBUFX3 U111 ( .A(n132), .Y(n114) );
  CLKBUFX3 U112 ( .A(n133), .Y(n113) );
  CLKBUFX3 U113 ( .A(n133), .Y(n112) );
  CLKBUFX3 U114 ( .A(n133), .Y(n111) );
  CLKBUFX3 U115 ( .A(n134), .Y(n110) );
  CLKBUFX3 U116 ( .A(n134), .Y(n109) );
  CLKBUFX3 U117 ( .A(n134), .Y(n108) );
  CLKBUFX3 U118 ( .A(n135), .Y(n107) );
  CLKBUFX3 U119 ( .A(n135), .Y(n106) );
  CLKBUFX3 U120 ( .A(n135), .Y(n105) );
  CLKBUFX3 U121 ( .A(n98), .Y(n97) );
  CLKBUFX3 U122 ( .A(n136), .Y(n104) );
  CLKBUFX3 U123 ( .A(n136), .Y(n103) );
  CLKBUFX3 U124 ( .A(n136), .Y(n102) );
  CLKBUFX3 U125 ( .A(n137), .Y(n101) );
  CLKBUFX3 U126 ( .A(n137), .Y(n100) );
  CLKBUFX3 U127 ( .A(n137), .Y(n99) );
  CLKBUFX3 U128 ( .A(n82), .Y(n128) );
  CLKBUFX3 U129 ( .A(n83), .Y(n129) );
  CLKBUFX3 U130 ( .A(n141), .Y(n130) );
  CLKBUFX3 U131 ( .A(n141), .Y(n131) );
  CLKBUFX3 U132 ( .A(n141), .Y(n132) );
  CLKBUFX3 U133 ( .A(n140), .Y(n133) );
  CLKBUFX3 U134 ( .A(n140), .Y(n134) );
  CLKBUFX3 U135 ( .A(n140), .Y(n135) );
  CLKBUFX3 U136 ( .A(n138), .Y(n98) );
  CLKBUFX3 U137 ( .A(n139), .Y(n138) );
  CLKBUFX3 U138 ( .A(n139), .Y(n136) );
  CLKBUFX3 U139 ( .A(n139), .Y(n137) );
  CLKBUFX3 U140 ( .A(n142), .Y(n141) );
  CLKBUFX3 U141 ( .A(n142), .Y(n140) );
  CLKBUFX3 U142 ( .A(n144), .Y(n142) );
  CLKBUFX3 U143 ( .A(n143), .Y(n139) );
  CLKBUFX3 U144 ( .A(n144), .Y(n143) );
  CLKBUFX3 U145 ( .A(clk), .Y(n144) );
  XOR2X1 U146 ( .A(out15[25]), .B(L14[25]), .Y(FP[25]) );
  XOR2X1 U147 ( .A(out15[17]), .B(L14[17]), .Y(FP[17]) );
  XOR2X1 U148 ( .A(out15[9]), .B(L14[9]), .Y(FP[9]) );
  XOR2X1 U149 ( .A(out15[1]), .B(L14[1]), .Y(FP[1]) );
  XOR2X1 U150 ( .A(out15[26]), .B(L14[26]), .Y(FP[26]) );
  XOR2X1 U151 ( .A(out15[18]), .B(L14[18]), .Y(FP[18]) );
  XOR2X1 U152 ( .A(out15[10]), .B(L14[10]), .Y(FP[10]) );
  XOR2X1 U153 ( .A(out15[2]), .B(L14[2]), .Y(FP[2]) );
  XOR2X1 U154 ( .A(out15[27]), .B(L14[27]), .Y(FP[27]) );
  XOR2X1 U155 ( .A(out15[19]), .B(L14[19]), .Y(FP[19]) );
  XOR2X1 U156 ( .A(out15[11]), .B(L14[11]), .Y(FP[11]) );
  XOR2X1 U157 ( .A(out15[3]), .B(L14[3]), .Y(FP[3]) );
  XOR2X1 U158 ( .A(out15[28]), .B(L14[28]), .Y(FP[28]) );
  XOR2X1 U159 ( .A(out15[20]), .B(L14[20]), .Y(FP[20]) );
  XOR2X1 U160 ( .A(out15[12]), .B(L14[12]), .Y(FP[12]) );
  XOR2X1 U161 ( .A(out15[4]), .B(L14[4]), .Y(FP[4]) );
  XOR2X1 U162 ( .A(out15[29]), .B(L14[29]), .Y(FP[29]) );
  XOR2X1 U163 ( .A(out15[21]), .B(L14[21]), .Y(FP[21]) );
  XOR2X1 U164 ( .A(out15[13]), .B(L14[13]), .Y(FP[13]) );
  XOR2X1 U165 ( .A(out15[5]), .B(L14[5]), .Y(FP[5]) );
  XOR2X1 U166 ( .A(out15[30]), .B(L14[30]), .Y(FP[30]) );
  XOR2X1 U167 ( .A(out15[22]), .B(L14[22]), .Y(FP[22]) );
  XOR2X1 U168 ( .A(out15[14]), .B(L14[14]), .Y(FP[14]) );
  XOR2X1 U169 ( .A(out15[6]), .B(L14[6]), .Y(FP[6]) );
  XOR2X1 U170 ( .A(out15[31]), .B(L14[31]), .Y(FP[31]) );
  XOR2X1 U171 ( .A(out15[23]), .B(L14[23]), .Y(FP[23]) );
  XOR2X1 U172 ( .A(out15[15]), .B(L14[15]), .Y(FP[15]) );
  XOR2X1 U173 ( .A(out15[7]), .B(L14[7]), .Y(FP[7]) );
  XOR2X1 U174 ( .A(out15[32]), .B(L14[32]), .Y(FP[32]) );
  XOR2X1 U175 ( .A(out15[24]), .B(L14[24]), .Y(FP[24]) );
  XOR2X1 U176 ( .A(out15[16]), .B(L14[16]), .Y(FP[16]) );
  XOR2X1 U177 ( .A(out15[8]), .B(L14[8]), .Y(FP[8]) );
  XOR2X1 U178 ( .A(out14[32]), .B(L13[32]), .Y(N479) );
  XOR2X1 U179 ( .A(out14[31]), .B(L13[31]), .Y(N478) );
  XOR2X1 U180 ( .A(out14[30]), .B(L13[30]), .Y(N477) );
  XOR2X1 U181 ( .A(out14[29]), .B(L13[29]), .Y(N476) );
  XOR2X1 U182 ( .A(out14[28]), .B(L13[28]), .Y(N475) );
  XOR2X1 U183 ( .A(out14[27]), .B(L13[27]), .Y(N474) );
  XOR2X1 U184 ( .A(out14[26]), .B(L13[26]), .Y(N473) );
  XOR2X1 U185 ( .A(out14[25]), .B(L13[25]), .Y(N472) );
  XOR2X1 U186 ( .A(out14[24]), .B(L13[24]), .Y(N471) );
  XOR2X1 U187 ( .A(out14[23]), .B(L13[23]), .Y(N470) );
  XOR2X1 U188 ( .A(out14[22]), .B(L13[22]), .Y(N469) );
  XOR2X1 U189 ( .A(out14[21]), .B(L13[21]), .Y(N468) );
  XOR2X1 U190 ( .A(out14[20]), .B(L13[20]), .Y(N467) );
  XOR2X1 U191 ( .A(out14[19]), .B(L13[19]), .Y(N466) );
  XOR2X1 U192 ( .A(out14[18]), .B(L13[18]), .Y(N465) );
  XOR2X1 U193 ( .A(out14[17]), .B(L13[17]), .Y(N464) );
  XOR2X1 U194 ( .A(out14[16]), .B(L13[16]), .Y(N463) );
  XOR2X1 U195 ( .A(out14[15]), .B(L13[15]), .Y(N462) );
  XOR2X1 U196 ( .A(out14[14]), .B(L13[14]), .Y(N461) );
  XOR2X1 U197 ( .A(out14[13]), .B(L13[13]), .Y(N460) );
  XOR2X1 U198 ( .A(out14[12]), .B(L13[12]), .Y(N459) );
  XOR2X1 U199 ( .A(out14[11]), .B(L13[11]), .Y(N458) );
  XOR2X1 U200 ( .A(out14[10]), .B(L13[10]), .Y(N457) );
  XOR2X1 U201 ( .A(out14[9]), .B(L13[9]), .Y(N456) );
  XOR2X1 U202 ( .A(out14[8]), .B(L13[8]), .Y(N455) );
  XOR2X1 U203 ( .A(out14[7]), .B(L13[7]), .Y(N454) );
  XOR2X1 U204 ( .A(out14[6]), .B(L13[6]), .Y(N453) );
  XOR2X1 U205 ( .A(out14[5]), .B(L13[5]), .Y(N452) );
  XOR2X1 U206 ( .A(out14[4]), .B(L13[4]), .Y(N451) );
  XOR2X1 U207 ( .A(out14[3]), .B(L13[3]), .Y(N450) );
  XOR2X1 U208 ( .A(out14[2]), .B(L13[2]), .Y(N449) );
  XOR2X1 U209 ( .A(out14[1]), .B(L13[1]), .Y(N448) );
  XOR2X1 U210 ( .A(out13[32]), .B(L12[32]), .Y(N447) );
  XOR2X1 U211 ( .A(out13[31]), .B(L12[31]), .Y(N446) );
  XOR2X1 U212 ( .A(out13[30]), .B(L12[30]), .Y(N445) );
  XOR2X1 U213 ( .A(out13[29]), .B(L12[29]), .Y(N444) );
  XOR2X1 U214 ( .A(out13[28]), .B(L12[28]), .Y(N443) );
  XOR2X1 U215 ( .A(out13[27]), .B(L12[27]), .Y(N442) );
  XOR2X1 U216 ( .A(out13[26]), .B(L12[26]), .Y(N441) );
  XOR2X1 U217 ( .A(out13[25]), .B(L12[25]), .Y(N440) );
  XOR2X1 U218 ( .A(out13[24]), .B(L12[24]), .Y(N439) );
  XOR2X1 U219 ( .A(out13[23]), .B(L12[23]), .Y(N438) );
  XOR2X1 U220 ( .A(out13[22]), .B(L12[22]), .Y(N437) );
  XOR2X1 U221 ( .A(out13[21]), .B(L12[21]), .Y(N436) );
  XOR2X1 U222 ( .A(out13[20]), .B(L12[20]), .Y(N435) );
  XOR2X1 U223 ( .A(out13[19]), .B(L12[19]), .Y(N434) );
  XOR2X1 U224 ( .A(out13[18]), .B(L12[18]), .Y(N433) );
  XOR2X1 U225 ( .A(out13[17]), .B(L12[17]), .Y(N432) );
  XOR2X1 U226 ( .A(out13[16]), .B(L12[16]), .Y(N431) );
  XOR2X1 U227 ( .A(out13[15]), .B(L12[15]), .Y(N430) );
  XOR2X1 U228 ( .A(out13[14]), .B(L12[14]), .Y(N429) );
  XOR2X1 U229 ( .A(out13[13]), .B(L12[13]), .Y(N428) );
  XOR2X1 U230 ( .A(out13[12]), .B(L12[12]), .Y(N427) );
  XOR2X1 U231 ( .A(out13[11]), .B(L12[11]), .Y(N426) );
  XOR2X1 U232 ( .A(out13[10]), .B(L12[10]), .Y(N425) );
  XOR2X1 U233 ( .A(out13[9]), .B(L12[9]), .Y(N424) );
  XOR2X1 U234 ( .A(out13[8]), .B(L12[8]), .Y(N423) );
  XOR2X1 U235 ( .A(out13[7]), .B(L12[7]), .Y(N422) );
  XOR2X1 U236 ( .A(out13[6]), .B(L12[6]), .Y(N421) );
  XOR2X1 U237 ( .A(out13[5]), .B(L12[5]), .Y(N420) );
  XOR2X1 U238 ( .A(out13[4]), .B(L12[4]), .Y(N419) );
  XOR2X1 U239 ( .A(out13[3]), .B(L12[3]), .Y(N418) );
  XOR2X1 U240 ( .A(out13[2]), .B(L12[2]), .Y(N417) );
  XOR2X1 U241 ( .A(out13[1]), .B(L12[1]), .Y(N416) );
  XOR2X1 U242 ( .A(out12[32]), .B(L11[32]), .Y(N415) );
  XOR2X1 U243 ( .A(out12[31]), .B(L11[31]), .Y(N414) );
  XOR2X1 U244 ( .A(out12[30]), .B(L11[30]), .Y(N413) );
  XOR2X1 U245 ( .A(out12[29]), .B(L11[29]), .Y(N412) );
  XOR2X1 U246 ( .A(out12[28]), .B(L11[28]), .Y(N411) );
  XOR2X1 U247 ( .A(out12[27]), .B(L11[27]), .Y(N410) );
  XOR2X1 U248 ( .A(out12[26]), .B(L11[26]), .Y(N409) );
  XOR2X1 U249 ( .A(out12[25]), .B(L11[25]), .Y(N408) );
  XOR2X1 U250 ( .A(out12[24]), .B(L11[24]), .Y(N407) );
  XOR2X1 U251 ( .A(out12[23]), .B(L11[23]), .Y(N406) );
  XOR2X1 U252 ( .A(out12[22]), .B(L11[22]), .Y(N405) );
  XOR2X1 U253 ( .A(out12[21]), .B(L11[21]), .Y(N404) );
  XOR2X1 U254 ( .A(out12[20]), .B(L11[20]), .Y(N403) );
  XOR2X1 U255 ( .A(out12[19]), .B(L11[19]), .Y(N402) );
  XOR2X1 U256 ( .A(out12[18]), .B(L11[18]), .Y(N401) );
  XOR2X1 U257 ( .A(out12[17]), .B(L11[17]), .Y(N400) );
  XOR2X1 U258 ( .A(out12[16]), .B(L11[16]), .Y(N399) );
  XOR2X1 U259 ( .A(out12[15]), .B(L11[15]), .Y(N398) );
  XOR2X1 U260 ( .A(out12[14]), .B(L11[14]), .Y(N397) );
  XOR2X1 U261 ( .A(out12[13]), .B(L11[13]), .Y(N396) );
  XOR2X1 U262 ( .A(out12[12]), .B(L11[12]), .Y(N395) );
  XOR2X1 U263 ( .A(out12[11]), .B(L11[11]), .Y(N394) );
  XOR2X1 U264 ( .A(out12[10]), .B(L11[10]), .Y(N393) );
  XOR2X1 U265 ( .A(out12[9]), .B(L11[9]), .Y(N392) );
  XOR2X1 U266 ( .A(out12[8]), .B(L11[8]), .Y(N391) );
  XOR2X1 U267 ( .A(out12[7]), .B(L11[7]), .Y(N390) );
  XOR2X1 U268 ( .A(out12[6]), .B(L11[6]), .Y(N389) );
  XOR2X1 U269 ( .A(out12[5]), .B(L11[5]), .Y(N388) );
  XOR2X1 U270 ( .A(out12[4]), .B(L11[4]), .Y(N387) );
  XOR2X1 U271 ( .A(out12[3]), .B(L11[3]), .Y(N386) );
  XOR2X1 U272 ( .A(out12[2]), .B(L11[2]), .Y(N385) );
  XOR2X1 U273 ( .A(out12[1]), .B(L11[1]), .Y(N384) );
  XOR2X1 U274 ( .A(out11[32]), .B(L10[32]), .Y(N383) );
  XOR2X1 U275 ( .A(out11[31]), .B(L10[31]), .Y(N382) );
  XOR2X1 U276 ( .A(out11[30]), .B(L10[30]), .Y(N381) );
  XOR2X1 U277 ( .A(out11[29]), .B(L10[29]), .Y(N380) );
  XOR2X1 U278 ( .A(out11[28]), .B(L10[28]), .Y(N379) );
  XOR2X1 U279 ( .A(out11[27]), .B(L10[27]), .Y(N378) );
  XOR2X1 U280 ( .A(out11[26]), .B(L10[26]), .Y(N377) );
  XOR2X1 U281 ( .A(out11[25]), .B(L10[25]), .Y(N376) );
  XOR2X1 U282 ( .A(out11[24]), .B(L10[24]), .Y(N375) );
  XOR2X1 U283 ( .A(out11[23]), .B(L10[23]), .Y(N374) );
  XOR2X1 U284 ( .A(out11[22]), .B(L10[22]), .Y(N373) );
  XOR2X1 U285 ( .A(out11[21]), .B(L10[21]), .Y(N372) );
  XOR2X1 U286 ( .A(out11[20]), .B(L10[20]), .Y(N371) );
  XOR2X1 U287 ( .A(out11[19]), .B(L10[19]), .Y(N370) );
  XOR2X1 U288 ( .A(out11[18]), .B(L10[18]), .Y(N369) );
  XOR2X1 U289 ( .A(out11[17]), .B(L10[17]), .Y(N368) );
  XOR2X1 U290 ( .A(out11[16]), .B(L10[16]), .Y(N367) );
  XOR2X1 U291 ( .A(out11[15]), .B(L10[15]), .Y(N366) );
  XOR2X1 U292 ( .A(out11[14]), .B(L10[14]), .Y(N365) );
  XOR2X1 U293 ( .A(out11[13]), .B(L10[13]), .Y(N364) );
  XOR2X1 U294 ( .A(out11[12]), .B(L10[12]), .Y(N363) );
  XOR2X1 U295 ( .A(out11[11]), .B(L10[11]), .Y(N362) );
  XOR2X1 U296 ( .A(out11[10]), .B(L10[10]), .Y(N361) );
  XOR2X1 U297 ( .A(out11[9]), .B(L10[9]), .Y(N360) );
  XOR2X1 U298 ( .A(out11[8]), .B(L10[8]), .Y(N359) );
  XOR2X1 U299 ( .A(out11[7]), .B(L10[7]), .Y(N358) );
  XOR2X1 U300 ( .A(out11[6]), .B(L10[6]), .Y(N357) );
  XOR2X1 U301 ( .A(out11[5]), .B(L10[5]), .Y(N356) );
  XOR2X1 U302 ( .A(out11[4]), .B(L10[4]), .Y(N355) );
  XOR2X1 U303 ( .A(out11[3]), .B(L10[3]), .Y(N354) );
  XOR2X1 U304 ( .A(out11[2]), .B(L10[2]), .Y(N353) );
  XOR2X1 U305 ( .A(out11[1]), .B(L10[1]), .Y(N352) );
  XOR2X1 U306 ( .A(out10[32]), .B(L9[32]), .Y(N351) );
  XOR2X1 U307 ( .A(out10[31]), .B(L9[31]), .Y(N350) );
  XOR2X1 U308 ( .A(out10[30]), .B(L9[30]), .Y(N349) );
  XOR2X1 U309 ( .A(out10[29]), .B(L9[29]), .Y(N348) );
  XOR2X1 U310 ( .A(out10[28]), .B(L9[28]), .Y(N347) );
  XOR2X1 U311 ( .A(out10[27]), .B(L9[27]), .Y(N346) );
  XOR2X1 U312 ( .A(out10[26]), .B(L9[26]), .Y(N345) );
  XOR2X1 U313 ( .A(out10[25]), .B(L9[25]), .Y(N344) );
  XOR2X1 U314 ( .A(out10[24]), .B(L9[24]), .Y(N343) );
  XOR2X1 U315 ( .A(out10[23]), .B(L9[23]), .Y(N342) );
  XOR2X1 U316 ( .A(out10[22]), .B(L9[22]), .Y(N341) );
  XOR2X1 U317 ( .A(out10[21]), .B(L9[21]), .Y(N340) );
  XOR2X1 U318 ( .A(out10[20]), .B(L9[20]), .Y(N339) );
  XOR2X1 U319 ( .A(out10[19]), .B(L9[19]), .Y(N338) );
  XOR2X1 U320 ( .A(out10[18]), .B(L9[18]), .Y(N337) );
  XOR2X1 U321 ( .A(out10[17]), .B(L9[17]), .Y(N336) );
  XOR2X1 U322 ( .A(out10[16]), .B(L9[16]), .Y(N335) );
  XOR2X1 U323 ( .A(out10[15]), .B(L9[15]), .Y(N334) );
  XOR2X1 U324 ( .A(out10[14]), .B(L9[14]), .Y(N333) );
  XOR2X1 U325 ( .A(out10[13]), .B(L9[13]), .Y(N332) );
  XOR2X1 U326 ( .A(out10[12]), .B(L9[12]), .Y(N331) );
  XOR2X1 U327 ( .A(out10[11]), .B(L9[11]), .Y(N330) );
  XOR2X1 U328 ( .A(out10[10]), .B(L9[10]), .Y(N329) );
  XOR2X1 U329 ( .A(out10[9]), .B(L9[9]), .Y(N328) );
  XOR2X1 U330 ( .A(out10[8]), .B(L9[8]), .Y(N327) );
  XOR2X1 U331 ( .A(out10[7]), .B(L9[7]), .Y(N326) );
  XOR2X1 U332 ( .A(out10[6]), .B(L9[6]), .Y(N325) );
  XOR2X1 U333 ( .A(out10[5]), .B(L9[5]), .Y(N324) );
  XOR2X1 U334 ( .A(out10[4]), .B(L9[4]), .Y(N323) );
  XOR2X1 U335 ( .A(out10[3]), .B(L9[3]), .Y(N322) );
  XOR2X1 U336 ( .A(out10[2]), .B(L9[2]), .Y(N321) );
  XOR2X1 U337 ( .A(out10[1]), .B(L9[1]), .Y(N320) );
  XOR2X1 U338 ( .A(out9[32]), .B(L8[32]), .Y(N319) );
  XOR2X1 U339 ( .A(out9[31]), .B(L8[31]), .Y(N318) );
  XOR2X1 U340 ( .A(out9[30]), .B(L8[30]), .Y(N317) );
  XOR2X1 U341 ( .A(out9[29]), .B(L8[29]), .Y(N316) );
  XOR2X1 U342 ( .A(out9[28]), .B(L8[28]), .Y(N315) );
  XOR2X1 U343 ( .A(out9[27]), .B(L8[27]), .Y(N314) );
  XOR2X1 U344 ( .A(out9[26]), .B(L8[26]), .Y(N313) );
  XOR2X1 U345 ( .A(out9[25]), .B(L8[25]), .Y(N312) );
  XOR2X1 U346 ( .A(out9[24]), .B(L8[24]), .Y(N311) );
  XOR2X1 U347 ( .A(out9[23]), .B(L8[23]), .Y(N310) );
  XOR2X1 U348 ( .A(out9[22]), .B(L8[22]), .Y(N309) );
  XOR2X1 U349 ( .A(out9[21]), .B(L8[21]), .Y(N308) );
  XOR2X1 U350 ( .A(out9[20]), .B(L8[20]), .Y(N307) );
  XOR2X1 U351 ( .A(out9[19]), .B(L8[19]), .Y(N306) );
  XOR2X1 U352 ( .A(out9[18]), .B(L8[18]), .Y(N305) );
  XOR2X1 U353 ( .A(out9[17]), .B(L8[17]), .Y(N304) );
  XOR2X1 U354 ( .A(out9[16]), .B(L8[16]), .Y(N303) );
  XOR2X1 U355 ( .A(out9[15]), .B(L8[15]), .Y(N302) );
  XOR2X1 U356 ( .A(out9[14]), .B(L8[14]), .Y(N301) );
  XOR2X1 U357 ( .A(out9[13]), .B(L8[13]), .Y(N300) );
  XOR2X1 U358 ( .A(out9[12]), .B(L8[12]), .Y(N299) );
  XOR2X1 U359 ( .A(out9[11]), .B(L8[11]), .Y(N298) );
  XOR2X1 U360 ( .A(out9[10]), .B(L8[10]), .Y(N297) );
  XOR2X1 U361 ( .A(out9[9]), .B(L8[9]), .Y(N296) );
  XOR2X1 U362 ( .A(out9[8]), .B(L8[8]), .Y(N295) );
  XOR2X1 U363 ( .A(out9[7]), .B(L8[7]), .Y(N294) );
  XOR2X1 U364 ( .A(out9[6]), .B(L8[6]), .Y(N293) );
  XOR2X1 U365 ( .A(out9[5]), .B(L8[5]), .Y(N292) );
  XOR2X1 U366 ( .A(out9[4]), .B(L8[4]), .Y(N291) );
  XOR2X1 U367 ( .A(out9[3]), .B(L8[3]), .Y(N290) );
  XOR2X1 U368 ( .A(out9[2]), .B(L8[2]), .Y(N289) );
  XOR2X1 U369 ( .A(out9[1]), .B(L8[1]), .Y(N288) );
  XOR2X1 U370 ( .A(out8[32]), .B(L7[32]), .Y(N287) );
  XOR2X1 U371 ( .A(out8[31]), .B(L7[31]), .Y(N286) );
  XOR2X1 U372 ( .A(out8[30]), .B(L7[30]), .Y(N285) );
  XOR2X1 U373 ( .A(out8[29]), .B(L7[29]), .Y(N284) );
  XOR2X1 U374 ( .A(out8[28]), .B(L7[28]), .Y(N283) );
  XOR2X1 U375 ( .A(out8[27]), .B(L7[27]), .Y(N282) );
  XOR2X1 U376 ( .A(out8[26]), .B(L7[26]), .Y(N281) );
  XOR2X1 U377 ( .A(out8[25]), .B(L7[25]), .Y(N280) );
  XOR2X1 U378 ( .A(out8[24]), .B(L7[24]), .Y(N279) );
  XOR2X1 U379 ( .A(out8[23]), .B(L7[23]), .Y(N278) );
  XOR2X1 U380 ( .A(out8[22]), .B(L7[22]), .Y(N277) );
  XOR2X1 U381 ( .A(out8[21]), .B(L7[21]), .Y(N276) );
  XOR2X1 U382 ( .A(out8[20]), .B(L7[20]), .Y(N275) );
  XOR2X1 U383 ( .A(out8[19]), .B(L7[19]), .Y(N274) );
  XOR2X1 U384 ( .A(out8[18]), .B(L7[18]), .Y(N273) );
  XOR2X1 U385 ( .A(out8[17]), .B(L7[17]), .Y(N272) );
  XOR2X1 U386 ( .A(out8[16]), .B(L7[16]), .Y(N271) );
  XOR2X1 U387 ( .A(out8[15]), .B(L7[15]), .Y(N270) );
  XOR2X1 U388 ( .A(out8[14]), .B(L7[14]), .Y(N269) );
  XOR2X1 U389 ( .A(out8[13]), .B(L7[13]), .Y(N268) );
  XOR2X1 U390 ( .A(out8[12]), .B(L7[12]), .Y(N267) );
  XOR2X1 U391 ( .A(out8[11]), .B(L7[11]), .Y(N266) );
  XOR2X1 U392 ( .A(out8[10]), .B(L7[10]), .Y(N265) );
  XOR2X1 U393 ( .A(out8[9]), .B(L7[9]), .Y(N264) );
  XOR2X1 U394 ( .A(out8[8]), .B(L7[8]), .Y(N263) );
  XOR2X1 U395 ( .A(out8[7]), .B(L7[7]), .Y(N262) );
  XOR2X1 U396 ( .A(out8[6]), .B(L7[6]), .Y(N261) );
  XOR2X1 U397 ( .A(out8[5]), .B(L7[5]), .Y(N260) );
  XOR2X1 U398 ( .A(out8[4]), .B(L7[4]), .Y(N259) );
  XOR2X1 U399 ( .A(out8[3]), .B(L7[3]), .Y(N258) );
  XOR2X1 U400 ( .A(out8[2]), .B(L7[2]), .Y(N257) );
  XOR2X1 U401 ( .A(out8[1]), .B(L7[1]), .Y(N256) );
  XOR2X1 U402 ( .A(out7[32]), .B(L6[32]), .Y(N255) );
  XOR2X1 U403 ( .A(out7[31]), .B(L6[31]), .Y(N254) );
  XOR2X1 U404 ( .A(out7[30]), .B(L6[30]), .Y(N253) );
  XOR2X1 U405 ( .A(out7[29]), .B(L6[29]), .Y(N252) );
  XOR2X1 U406 ( .A(out7[28]), .B(L6[28]), .Y(N251) );
  XOR2X1 U407 ( .A(out7[27]), .B(L6[27]), .Y(N250) );
  XOR2X1 U408 ( .A(out7[26]), .B(L6[26]), .Y(N249) );
  XOR2X1 U409 ( .A(out7[25]), .B(L6[25]), .Y(N248) );
  XOR2X1 U410 ( .A(out7[24]), .B(L6[24]), .Y(N247) );
  XOR2X1 U411 ( .A(out7[23]), .B(L6[23]), .Y(N246) );
  XOR2X1 U412 ( .A(out7[22]), .B(L6[22]), .Y(N245) );
  XOR2X1 U413 ( .A(out7[21]), .B(L6[21]), .Y(N244) );
  XOR2X1 U414 ( .A(out7[20]), .B(L6[20]), .Y(N243) );
  XOR2X1 U415 ( .A(out7[19]), .B(L6[19]), .Y(N242) );
  XOR2X1 U416 ( .A(out7[18]), .B(L6[18]), .Y(N241) );
  XOR2X1 U417 ( .A(out7[17]), .B(L6[17]), .Y(N240) );
  XOR2X1 U418 ( .A(out7[16]), .B(L6[16]), .Y(N239) );
  XOR2X1 U419 ( .A(out7[15]), .B(L6[15]), .Y(N238) );
  XOR2X1 U420 ( .A(out7[14]), .B(L6[14]), .Y(N237) );
  XOR2X1 U421 ( .A(out7[13]), .B(L6[13]), .Y(N236) );
  XOR2X1 U422 ( .A(out7[12]), .B(L6[12]), .Y(N235) );
  XOR2X1 U423 ( .A(out7[11]), .B(L6[11]), .Y(N234) );
  XOR2X1 U424 ( .A(out7[10]), .B(L6[10]), .Y(N233) );
  XOR2X1 U425 ( .A(out7[9]), .B(L6[9]), .Y(N232) );
  XOR2X1 U426 ( .A(out7[8]), .B(L6[8]), .Y(N231) );
  XOR2X1 U427 ( .A(out7[7]), .B(L6[7]), .Y(N230) );
  XOR2X1 U428 ( .A(out7[6]), .B(L6[6]), .Y(N229) );
  XOR2X1 U429 ( .A(out7[5]), .B(L6[5]), .Y(N228) );
  XOR2X1 U430 ( .A(out7[4]), .B(L6[4]), .Y(N227) );
  XOR2X1 U431 ( .A(out7[3]), .B(L6[3]), .Y(N226) );
  XOR2X1 U432 ( .A(out7[2]), .B(L6[2]), .Y(N225) );
  XOR2X1 U433 ( .A(out7[1]), .B(L6[1]), .Y(N224) );
  XOR2X1 U434 ( .A(out6[32]), .B(L5[32]), .Y(N223) );
  XOR2X1 U435 ( .A(out6[31]), .B(L5[31]), .Y(N222) );
  XOR2X1 U436 ( .A(out6[30]), .B(L5[30]), .Y(N221) );
  XOR2X1 U437 ( .A(out6[29]), .B(L5[29]), .Y(N220) );
  XOR2X1 U438 ( .A(out6[28]), .B(L5[28]), .Y(N219) );
  XOR2X1 U439 ( .A(out6[27]), .B(L5[27]), .Y(N218) );
  XOR2X1 U440 ( .A(out6[26]), .B(L5[26]), .Y(N217) );
  XOR2X1 U441 ( .A(out6[25]), .B(L5[25]), .Y(N216) );
  XOR2X1 U442 ( .A(out6[24]), .B(L5[24]), .Y(N215) );
  XOR2X1 U443 ( .A(out6[23]), .B(L5[23]), .Y(N214) );
  XOR2X1 U444 ( .A(out6[22]), .B(L5[22]), .Y(N213) );
  XOR2X1 U445 ( .A(out6[21]), .B(L5[21]), .Y(N212) );
  XOR2X1 U446 ( .A(out6[20]), .B(L5[20]), .Y(N211) );
  XOR2X1 U447 ( .A(out6[19]), .B(L5[19]), .Y(N210) );
  XOR2X1 U448 ( .A(out6[18]), .B(L5[18]), .Y(N209) );
  XOR2X1 U449 ( .A(out6[17]), .B(L5[17]), .Y(N208) );
  XOR2X1 U450 ( .A(out6[16]), .B(L5[16]), .Y(N207) );
  XOR2X1 U451 ( .A(out6[15]), .B(L5[15]), .Y(N206) );
  XOR2X1 U452 ( .A(out6[14]), .B(L5[14]), .Y(N205) );
  XOR2X1 U453 ( .A(out6[13]), .B(L5[13]), .Y(N204) );
  XOR2X1 U454 ( .A(out6[12]), .B(L5[12]), .Y(N203) );
  XOR2X1 U455 ( .A(out6[11]), .B(L5[11]), .Y(N202) );
  XOR2X1 U456 ( .A(out6[10]), .B(L5[10]), .Y(N201) );
  XOR2X1 U457 ( .A(out6[9]), .B(L5[9]), .Y(N200) );
  XOR2X1 U458 ( .A(out6[8]), .B(L5[8]), .Y(N199) );
  XOR2X1 U459 ( .A(out6[7]), .B(L5[7]), .Y(N198) );
  XOR2X1 U460 ( .A(out6[6]), .B(L5[6]), .Y(N197) );
  XOR2X1 U461 ( .A(out6[5]), .B(L5[5]), .Y(N196) );
  XOR2X1 U462 ( .A(out6[4]), .B(L5[4]), .Y(N195) );
  XOR2X1 U463 ( .A(out6[3]), .B(L5[3]), .Y(N194) );
  XOR2X1 U464 ( .A(out6[2]), .B(L5[2]), .Y(N193) );
  XOR2X1 U465 ( .A(out6[1]), .B(L5[1]), .Y(N192) );
  XOR2X1 U466 ( .A(out5[32]), .B(L4[32]), .Y(N191) );
  XOR2X1 U467 ( .A(out5[31]), .B(L4[31]), .Y(N190) );
  XOR2X1 U468 ( .A(out5[30]), .B(L4[30]), .Y(N189) );
  XOR2X1 U469 ( .A(out5[29]), .B(L4[29]), .Y(N188) );
  XOR2X1 U470 ( .A(out5[28]), .B(L4[28]), .Y(N187) );
  XOR2X1 U471 ( .A(out5[27]), .B(L4[27]), .Y(N186) );
  XOR2X1 U472 ( .A(out5[26]), .B(L4[26]), .Y(N185) );
  XOR2X1 U473 ( .A(out5[25]), .B(L4[25]), .Y(N184) );
  XOR2X1 U474 ( .A(out5[24]), .B(L4[24]), .Y(N183) );
  XOR2X1 U475 ( .A(out5[23]), .B(L4[23]), .Y(N182) );
  XOR2X1 U476 ( .A(out5[22]), .B(L4[22]), .Y(N181) );
  XOR2X1 U477 ( .A(out5[21]), .B(L4[21]), .Y(N180) );
  XOR2X1 U478 ( .A(out5[20]), .B(L4[20]), .Y(N179) );
  XOR2X1 U479 ( .A(out5[19]), .B(L4[19]), .Y(N178) );
  XOR2X1 U480 ( .A(out5[18]), .B(L4[18]), .Y(N177) );
  XOR2X1 U481 ( .A(out5[17]), .B(L4[17]), .Y(N176) );
  XOR2X1 U482 ( .A(out5[16]), .B(L4[16]), .Y(N175) );
  XOR2X1 U483 ( .A(out5[15]), .B(L4[15]), .Y(N174) );
  XOR2X1 U484 ( .A(out5[14]), .B(L4[14]), .Y(N173) );
  XOR2X1 U485 ( .A(out5[13]), .B(L4[13]), .Y(N172) );
  XOR2X1 U486 ( .A(out5[12]), .B(L4[12]), .Y(N171) );
  XOR2X1 U487 ( .A(out5[11]), .B(L4[11]), .Y(N170) );
  XOR2X1 U488 ( .A(out5[10]), .B(L4[10]), .Y(N169) );
  XOR2X1 U489 ( .A(out5[9]), .B(L4[9]), .Y(N168) );
  XOR2X1 U490 ( .A(out5[8]), .B(L4[8]), .Y(N167) );
  XOR2X1 U491 ( .A(out5[7]), .B(L4[7]), .Y(N166) );
  XOR2X1 U492 ( .A(out5[6]), .B(L4[6]), .Y(N165) );
  XOR2X1 U493 ( .A(out5[5]), .B(L4[5]), .Y(N164) );
  XOR2X1 U494 ( .A(out5[4]), .B(L4[4]), .Y(N163) );
  XOR2X1 U495 ( .A(out5[3]), .B(L4[3]), .Y(N162) );
  XOR2X1 U496 ( .A(out5[2]), .B(L4[2]), .Y(N161) );
  XOR2X1 U497 ( .A(out5[1]), .B(L4[1]), .Y(N160) );
  XOR2X1 U498 ( .A(out4[32]), .B(L3[32]), .Y(N159) );
  XOR2X1 U499 ( .A(out4[31]), .B(L3[31]), .Y(N158) );
  XOR2X1 U500 ( .A(out4[30]), .B(L3[30]), .Y(N157) );
  XOR2X1 U501 ( .A(out4[29]), .B(L3[29]), .Y(N156) );
  XOR2X1 U502 ( .A(out4[28]), .B(L3[28]), .Y(N155) );
  XOR2X1 U503 ( .A(out4[27]), .B(L3[27]), .Y(N154) );
  XOR2X1 U504 ( .A(out4[26]), .B(L3[26]), .Y(N153) );
  XOR2X1 U505 ( .A(out4[25]), .B(L3[25]), .Y(N152) );
  XOR2X1 U506 ( .A(out4[24]), .B(L3[24]), .Y(N151) );
  XOR2X1 U507 ( .A(out4[23]), .B(L3[23]), .Y(N150) );
  XOR2X1 U508 ( .A(out4[22]), .B(L3[22]), .Y(N149) );
  XOR2X1 U509 ( .A(out4[21]), .B(L3[21]), .Y(N148) );
  XOR2X1 U510 ( .A(out4[20]), .B(L3[20]), .Y(N147) );
  XOR2X1 U511 ( .A(out4[19]), .B(L3[19]), .Y(N146) );
  XOR2X1 U512 ( .A(out4[18]), .B(L3[18]), .Y(N145) );
  XOR2X1 U513 ( .A(out4[17]), .B(L3[17]), .Y(N144) );
  XOR2X1 U514 ( .A(out4[16]), .B(L3[16]), .Y(N143) );
  XOR2X1 U515 ( .A(out4[15]), .B(L3[15]), .Y(N142) );
  XOR2X1 U516 ( .A(out4[14]), .B(L3[14]), .Y(N141) );
  XOR2X1 U517 ( .A(out4[13]), .B(L3[13]), .Y(N140) );
  XOR2X1 U518 ( .A(out4[12]), .B(L3[12]), .Y(N139) );
  XOR2X1 U519 ( .A(out4[11]), .B(L3[11]), .Y(N138) );
  XOR2X1 U520 ( .A(out4[10]), .B(L3[10]), .Y(N137) );
  XOR2X1 U521 ( .A(out4[9]), .B(L3[9]), .Y(N136) );
  XOR2X1 U522 ( .A(out4[8]), .B(L3[8]), .Y(N135) );
  XOR2X1 U523 ( .A(out4[7]), .B(L3[7]), .Y(N134) );
  XOR2X1 U524 ( .A(out4[6]), .B(L3[6]), .Y(N133) );
  XOR2X1 U525 ( .A(out4[5]), .B(L3[5]), .Y(N132) );
  XOR2X1 U526 ( .A(out4[4]), .B(L3[4]), .Y(N131) );
  XOR2X1 U527 ( .A(out4[3]), .B(L3[3]), .Y(N130) );
  XOR2X1 U528 ( .A(out4[2]), .B(L3[2]), .Y(N129) );
  XOR2X1 U529 ( .A(out4[1]), .B(L3[1]), .Y(N128) );
  XOR2X1 U530 ( .A(out3[32]), .B(L2[32]), .Y(N127) );
  XOR2X1 U531 ( .A(out3[31]), .B(L2[31]), .Y(N126) );
  XOR2X1 U532 ( .A(out3[30]), .B(L2[30]), .Y(N125) );
  XOR2X1 U533 ( .A(out3[29]), .B(L2[29]), .Y(N124) );
  XOR2X1 U534 ( .A(out3[28]), .B(L2[28]), .Y(N123) );
  XOR2X1 U535 ( .A(out3[27]), .B(L2[27]), .Y(N122) );
  XOR2X1 U536 ( .A(out3[26]), .B(L2[26]), .Y(N121) );
  XOR2X1 U537 ( .A(out3[25]), .B(L2[25]), .Y(N120) );
  XOR2X1 U538 ( .A(out3[24]), .B(L2[24]), .Y(N119) );
  XOR2X1 U539 ( .A(out3[23]), .B(L2[23]), .Y(N118) );
  XOR2X1 U540 ( .A(out3[22]), .B(L2[22]), .Y(N117) );
  XOR2X1 U541 ( .A(out3[21]), .B(L2[21]), .Y(N116) );
  XOR2X1 U542 ( .A(out3[20]), .B(L2[20]), .Y(N115) );
  XOR2X1 U543 ( .A(out3[19]), .B(L2[19]), .Y(N114) );
  XOR2X1 U544 ( .A(out3[18]), .B(L2[18]), .Y(N113) );
  XOR2X1 U545 ( .A(out3[17]), .B(L2[17]), .Y(N112) );
  XOR2X1 U546 ( .A(out3[16]), .B(L2[16]), .Y(N111) );
  XOR2X1 U547 ( .A(out3[15]), .B(L2[15]), .Y(N110) );
  XOR2X1 U548 ( .A(out3[14]), .B(L2[14]), .Y(N109) );
  XOR2X1 U549 ( .A(out3[13]), .B(L2[13]), .Y(N108) );
  XOR2X1 U550 ( .A(out3[12]), .B(L2[12]), .Y(N107) );
  XOR2X1 U551 ( .A(out3[11]), .B(L2[11]), .Y(N106) );
  XOR2X1 U552 ( .A(out3[10]), .B(L2[10]), .Y(N105) );
  XOR2X1 U553 ( .A(out3[9]), .B(L2[9]), .Y(N104) );
  XOR2X1 U554 ( .A(out3[8]), .B(L2[8]), .Y(N103) );
  XOR2X1 U555 ( .A(out3[7]), .B(L2[7]), .Y(N102) );
  XOR2X1 U556 ( .A(out3[6]), .B(L2[6]), .Y(N101) );
  XOR2X1 U557 ( .A(out3[5]), .B(L2[5]), .Y(N100) );
  XOR2X1 U558 ( .A(out3[4]), .B(L2[4]), .Y(N99) );
  XOR2X1 U559 ( .A(out3[3]), .B(L2[3]), .Y(N98) );
  XOR2X1 U560 ( .A(out3[2]), .B(L2[2]), .Y(N97) );
  XOR2X1 U561 ( .A(out3[1]), .B(L2[1]), .Y(N96) );
  XOR2X1 U562 ( .A(out2[32]), .B(L1[32]), .Y(N95) );
  XOR2X1 U563 ( .A(out2[31]), .B(L1[31]), .Y(N94) );
  XOR2X1 U564 ( .A(out2[30]), .B(L1[30]), .Y(N93) );
  XOR2X1 U565 ( .A(out2[29]), .B(L1[29]), .Y(N92) );
  XOR2X1 U566 ( .A(out2[28]), .B(L1[28]), .Y(N91) );
  XOR2X1 U567 ( .A(out2[27]), .B(L1[27]), .Y(N90) );
  XOR2X1 U568 ( .A(out2[26]), .B(L1[26]), .Y(N89) );
  XOR2X1 U569 ( .A(out2[25]), .B(L1[25]), .Y(N88) );
  XOR2X1 U570 ( .A(out2[24]), .B(L1[24]), .Y(N87) );
  XOR2X1 U571 ( .A(out2[23]), .B(L1[23]), .Y(N86) );
  XOR2X1 U572 ( .A(out2[22]), .B(L1[22]), .Y(N85) );
  XOR2X1 U573 ( .A(out2[21]), .B(L1[21]), .Y(N84) );
  XOR2X1 U574 ( .A(out2[20]), .B(L1[20]), .Y(N83) );
  XOR2X1 U575 ( .A(out2[19]), .B(L1[19]), .Y(N82) );
  XOR2X1 U576 ( .A(out2[18]), .B(L1[18]), .Y(N81) );
  XOR2X1 U577 ( .A(out2[17]), .B(L1[17]), .Y(N80) );
  XOR2X1 U578 ( .A(out2[16]), .B(L1[16]), .Y(N79) );
  XOR2X1 U579 ( .A(out2[15]), .B(L1[15]), .Y(N78) );
  XOR2X1 U580 ( .A(out2[14]), .B(L1[14]), .Y(N77) );
  XOR2X1 U581 ( .A(out2[13]), .B(L1[13]), .Y(N76) );
  XOR2X1 U582 ( .A(out2[12]), .B(L1[12]), .Y(N75) );
  XOR2X1 U583 ( .A(out2[11]), .B(L1[11]), .Y(N74) );
  XOR2X1 U584 ( .A(out2[10]), .B(L1[10]), .Y(N73) );
  XOR2X1 U585 ( .A(out2[9]), .B(L1[9]), .Y(N72) );
  XOR2X1 U586 ( .A(out2[8]), .B(L1[8]), .Y(N71) );
  XOR2X1 U587 ( .A(out2[7]), .B(L1[7]), .Y(N70) );
  XOR2X1 U588 ( .A(out2[6]), .B(L1[6]), .Y(N69) );
  XOR2X1 U589 ( .A(out2[5]), .B(L1[5]), .Y(N68) );
  XOR2X1 U590 ( .A(out2[4]), .B(L1[4]), .Y(N67) );
  XOR2X1 U591 ( .A(out2[3]), .B(L1[3]), .Y(N66) );
  XOR2X1 U592 ( .A(out2[2]), .B(L1[2]), .Y(N65) );
  XOR2X1 U593 ( .A(out2[1]), .B(L1[1]), .Y(N64) );
  XOR2X1 U594 ( .A(out1[32]), .B(L0[32]), .Y(N63) );
  XOR2X1 U595 ( .A(out1[31]), .B(L0[31]), .Y(N62) );
  XOR2X1 U596 ( .A(out1[30]), .B(L0[30]), .Y(N61) );
  XOR2X1 U597 ( .A(out1[29]), .B(L0[29]), .Y(N60) );
  XOR2X1 U598 ( .A(out1[28]), .B(L0[28]), .Y(N59) );
  XOR2X1 U599 ( .A(out1[27]), .B(L0[27]), .Y(N58) );
  XOR2X1 U600 ( .A(out1[26]), .B(L0[26]), .Y(N57) );
  XOR2X1 U601 ( .A(out1[25]), .B(L0[25]), .Y(N56) );
  XOR2X1 U602 ( .A(out1[24]), .B(L0[24]), .Y(N55) );
  XOR2X1 U603 ( .A(out1[23]), .B(L0[23]), .Y(N54) );
  XOR2X1 U604 ( .A(out1[22]), .B(L0[22]), .Y(N53) );
  XOR2X1 U605 ( .A(out1[21]), .B(L0[21]), .Y(N52) );
  XOR2X1 U606 ( .A(out1[20]), .B(L0[20]), .Y(N51) );
  XOR2X1 U607 ( .A(out1[19]), .B(L0[19]), .Y(N50) );
  XOR2X1 U608 ( .A(out1[18]), .B(L0[18]), .Y(N49) );
  XOR2X1 U609 ( .A(out1[17]), .B(L0[17]), .Y(N48) );
  XOR2X1 U610 ( .A(out1[16]), .B(L0[16]), .Y(N47) );
  XOR2X1 U611 ( .A(out1[15]), .B(L0[15]), .Y(N46) );
  XOR2X1 U612 ( .A(out1[14]), .B(L0[14]), .Y(N45) );
  XOR2X1 U613 ( .A(out1[13]), .B(L0[13]), .Y(N44) );
  XOR2X1 U614 ( .A(out1[12]), .B(L0[12]), .Y(N43) );
  XOR2X1 U615 ( .A(out1[11]), .B(L0[11]), .Y(N42) );
  XOR2X1 U616 ( .A(out1[10]), .B(L0[10]), .Y(N41) );
  XOR2X1 U617 ( .A(out1[9]), .B(L0[9]), .Y(N40) );
  XOR2X1 U618 ( .A(out1[8]), .B(L0[8]), .Y(N39) );
  XOR2X1 U619 ( .A(out1[7]), .B(L0[7]), .Y(N38) );
  XOR2X1 U620 ( .A(out1[6]), .B(L0[6]), .Y(N37) );
  XOR2X1 U621 ( .A(out1[5]), .B(L0[5]), .Y(N36) );
  XOR2X1 U622 ( .A(out1[4]), .B(L0[4]), .Y(N35) );
  XOR2X1 U623 ( .A(out1[3]), .B(L0[3]), .Y(N34) );
  XOR2X1 U624 ( .A(out1[2]), .B(L0[2]), .Y(N33) );
  XOR2X1 U625 ( .A(out1[1]), .B(L0[1]), .Y(N32) );
  XOR2X1 U626 ( .A(out0[32]), .B(desIn_r[56]), .Y(N31) );
  XOR2X1 U627 ( .A(out0[31]), .B(desIn_r[48]), .Y(N30) );
  XOR2X1 U628 ( .A(out0[30]), .B(desIn_r[40]), .Y(N29) );
  XOR2X1 U629 ( .A(out0[29]), .B(desIn_r[32]), .Y(N28) );
  XOR2X1 U630 ( .A(out0[28]), .B(desIn_r[24]), .Y(N27) );
  XOR2X1 U631 ( .A(out0[27]), .B(desIn_r[16]), .Y(N26) );
  XOR2X1 U632 ( .A(out0[26]), .B(desIn_r[8]), .Y(N25) );
  XOR2X1 U633 ( .A(out0[25]), .B(desIn_r[0]), .Y(N24) );
  XOR2X1 U634 ( .A(out0[24]), .B(desIn_r[58]), .Y(N23) );
  XOR2X1 U635 ( .A(out0[23]), .B(desIn_r[50]), .Y(N22) );
  XOR2X1 U636 ( .A(out0[22]), .B(desIn_r[42]), .Y(N21) );
  XOR2X1 U637 ( .A(out0[21]), .B(desIn_r[34]), .Y(N20) );
  XOR2X1 U638 ( .A(out0[20]), .B(desIn_r[26]), .Y(N19) );
  XOR2X1 U639 ( .A(out0[19]), .B(desIn_r[18]), .Y(N18) );
  XOR2X1 U640 ( .A(out0[18]), .B(desIn_r[10]), .Y(N17) );
  XOR2X1 U641 ( .A(out0[17]), .B(desIn_r[2]), .Y(N16) );
  XOR2X1 U642 ( .A(out0[16]), .B(desIn_r[60]), .Y(N15) );
  XOR2X1 U643 ( .A(out0[15]), .B(desIn_r[52]), .Y(N14) );
  XOR2X1 U644 ( .A(out0[14]), .B(desIn_r[44]), .Y(N13) );
  XOR2X1 U645 ( .A(out0[13]), .B(desIn_r[36]), .Y(N12) );
  XOR2X1 U646 ( .A(out0[12]), .B(desIn_r[28]), .Y(N11) );
  XOR2X1 U647 ( .A(out0[11]), .B(desIn_r[20]), .Y(N10) );
  XOR2X1 U648 ( .A(out0[10]), .B(desIn_r[12]), .Y(N9) );
  XOR2X1 U649 ( .A(out0[9]), .B(desIn_r[4]), .Y(N8) );
  XOR2X1 U650 ( .A(out0[8]), .B(desIn_r[62]), .Y(N7) );
  XOR2X1 U651 ( .A(out0[7]), .B(desIn_r[54]), .Y(N6) );
  XOR2X1 U652 ( .A(out0[6]), .B(desIn_r[46]), .Y(N5) );
  XOR2X1 U653 ( .A(out0[5]), .B(desIn_r[38]), .Y(N4) );
  XOR2X1 U654 ( .A(out0[4]), .B(desIn_r[30]), .Y(N3) );
  XOR2X1 U655 ( .A(out0[3]), .B(desIn_r[22]), .Y(N2) );
  XOR2X1 U656 ( .A(out0[2]), .B(desIn_r[14]), .Y(N1) );
  XOR2X1 U657 ( .A(out0[1]), .B(desIn_r[6]), .Y(N0) );
  CLKBUFX3 U658 ( .A(decrypt), .Y(n1) );
endmodule


module des2 ( desIn, key1, key2, decrypt, desEnable, reset_n, clk, desOut );
  input [63:0] desIn;
  input [55:0] key1;
  input [55:0] key2;
  output [63:0] desOut;
  input decrypt, desEnable, reset_n, clk;
  wire   N3, N6, N7, N8, N10, N11, N12, N13, N14, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         \add_24/carry[4] , \add_24/carry[3] , \add_24/carry[2] , n1, n2, n3,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330;
  wire   [4:0] cnt;
  wire   [63:0] din;
  wire   [55:0] key;

  des d2 ( .desOut(desOut), .desIn(din), .key(key), .decrypt(decrypt), .clk(
        n208) );
  ADDHX1 \add_24/U1_1_1  ( .A(cnt[1]), .B(cnt[0]), .CO(\add_24/carry[2] ), .S(
        N6) );
  ADDHX1 \add_24/U1_1_2  ( .A(cnt[2]), .B(\add_24/carry[2] ), .CO(
        \add_24/carry[3] ), .S(N7) );
  ADDHX1 \add_24/U1_1_3  ( .A(cnt[3]), .B(\add_24/carry[3] ), .CO(
        \add_24/carry[4] ), .S(N8) );
  DFFRX1 flag_reg ( .D(n127), .CK(n203), .RN(n138), .QN(n126) );
  DFFRX1 \cnt_reg[1]  ( .D(N11), .CK(n203), .RN(n138), .Q(cnt[1]) );
  DFFRX1 \cnt_reg[4]  ( .D(N14), .CK(n203), .RN(n138), .Q(cnt[4]), .QN(n2) );
  DFFRX1 \key_reg[55]  ( .D(n275), .CK(n203), .RN(n138), .Q(key[55]) );
  DFFRX1 \key_reg[54]  ( .D(n276), .CK(n202), .RN(n138), .Q(key[54]) );
  DFFRX1 \key_reg[53]  ( .D(n277), .CK(n202), .RN(n138), .Q(key[53]) );
  DFFRX1 \key_reg[52]  ( .D(n278), .CK(n202), .RN(n137), .Q(key[52]) );
  DFFRX1 \key_reg[51]  ( .D(n279), .CK(n202), .RN(n137), .Q(key[51]) );
  DFFRX1 \key_reg[50]  ( .D(n280), .CK(n202), .RN(n137), .Q(key[50]) );
  DFFRX1 \key_reg[49]  ( .D(n281), .CK(n202), .RN(n137), .Q(key[49]) );
  DFFRX1 \key_reg[48]  ( .D(n282), .CK(n202), .RN(n137), .Q(key[48]) );
  DFFRX1 \key_reg[47]  ( .D(n283), .CK(n202), .RN(n137), .Q(key[47]) );
  DFFRX1 \key_reg[46]  ( .D(n284), .CK(n202), .RN(n137), .Q(key[46]) );
  DFFRX1 \key_reg[45]  ( .D(n285), .CK(n202), .RN(n137), .Q(key[45]) );
  DFFRX1 \key_reg[44]  ( .D(n286), .CK(n201), .RN(n137), .Q(key[44]) );
  DFFRX1 \key_reg[43]  ( .D(n287), .CK(n201), .RN(n136), .Q(key[43]) );
  DFFRX1 \key_reg[42]  ( .D(n288), .CK(n201), .RN(n136), .Q(key[42]) );
  DFFRX1 \key_reg[41]  ( .D(n289), .CK(n201), .RN(n136), .Q(key[41]) );
  DFFRX1 \key_reg[40]  ( .D(n290), .CK(n201), .RN(n136), .Q(key[40]) );
  DFFRX1 \key_reg[39]  ( .D(n291), .CK(n201), .RN(n136), .Q(key[39]) );
  DFFRX1 \key_reg[38]  ( .D(n292), .CK(n201), .RN(n136), .Q(key[38]) );
  DFFRX1 \key_reg[37]  ( .D(n293), .CK(n201), .RN(n136), .Q(key[37]) );
  DFFRX1 \key_reg[36]  ( .D(n294), .CK(n201), .RN(n136), .Q(key[36]) );
  DFFRX1 \key_reg[35]  ( .D(n295), .CK(n201), .RN(n136), .Q(key[35]) );
  DFFRX1 \key_reg[34]  ( .D(n296), .CK(n200), .RN(n135), .Q(key[34]) );
  DFFRX1 \key_reg[33]  ( .D(n297), .CK(n200), .RN(n135), .Q(key[33]) );
  DFFRX1 \key_reg[32]  ( .D(n298), .CK(n200), .RN(n135), .Q(key[32]) );
  DFFRX1 \key_reg[31]  ( .D(n299), .CK(n200), .RN(n135), .Q(key[31]) );
  DFFRX1 \key_reg[30]  ( .D(n300), .CK(n200), .RN(n135), .Q(key[30]) );
  DFFRX1 \key_reg[29]  ( .D(n301), .CK(n200), .RN(n135), .Q(key[29]) );
  DFFRX1 \key_reg[28]  ( .D(n302), .CK(n200), .RN(n135), .Q(key[28]) );
  DFFRX1 \key_reg[27]  ( .D(n303), .CK(n200), .RN(n135), .Q(key[27]) );
  DFFRX1 \key_reg[26]  ( .D(n304), .CK(n200), .RN(n135), .Q(key[26]) );
  DFFRX1 \key_reg[25]  ( .D(n305), .CK(n200), .RN(n134), .Q(key[25]) );
  DFFRX1 \key_reg[24]  ( .D(n306), .CK(n199), .RN(n134), .Q(key[24]) );
  DFFRX1 \key_reg[23]  ( .D(n307), .CK(n199), .RN(n134), .Q(key[23]) );
  DFFRX1 \key_reg[22]  ( .D(n308), .CK(n199), .RN(n134), .Q(key[22]) );
  DFFRX1 \key_reg[21]  ( .D(n309), .CK(n199), .RN(n134), .Q(key[21]) );
  DFFRX1 \key_reg[20]  ( .D(n310), .CK(n199), .RN(n134), .Q(key[20]) );
  DFFRX1 \key_reg[19]  ( .D(n311), .CK(n199), .RN(n134), .Q(key[19]) );
  DFFRX1 \key_reg[18]  ( .D(n312), .CK(n199), .RN(n134), .Q(key[18]) );
  DFFRX1 \key_reg[17]  ( .D(n313), .CK(n199), .RN(n134), .Q(key[17]) );
  DFFRX1 \key_reg[16]  ( .D(n314), .CK(n199), .RN(n133), .Q(key[16]) );
  DFFRX1 \key_reg[15]  ( .D(n315), .CK(n199), .RN(n133), .Q(key[15]) );
  DFFRX1 \key_reg[14]  ( .D(n316), .CK(n198), .RN(n133), .Q(key[14]) );
  DFFRX1 \key_reg[13]  ( .D(n317), .CK(n198), .RN(n133), .Q(key[13]) );
  DFFRX1 \key_reg[12]  ( .D(n318), .CK(n198), .RN(n133), .Q(key[12]) );
  DFFRX1 \key_reg[11]  ( .D(n319), .CK(n198), .RN(n133), .Q(key[11]) );
  DFFRX1 \key_reg[10]  ( .D(n320), .CK(n198), .RN(n133), .Q(key[10]) );
  DFFRX1 \key_reg[9]  ( .D(n321), .CK(n198), .RN(n133), .Q(key[9]) );
  DFFRX1 \key_reg[8]  ( .D(n322), .CK(n198), .RN(n133), .Q(key[8]) );
  DFFRX1 \key_reg[7]  ( .D(n323), .CK(n198), .RN(n132), .Q(key[7]) );
  DFFRX1 \key_reg[6]  ( .D(n324), .CK(n198), .RN(n132), .Q(key[6]) );
  DFFRX1 \key_reg[5]  ( .D(n325), .CK(n198), .RN(n132), .Q(key[5]) );
  DFFRX1 \key_reg[4]  ( .D(n326), .CK(n197), .RN(n132), .Q(key[4]) );
  DFFRX1 \key_reg[3]  ( .D(n327), .CK(n197), .RN(n132), .Q(key[3]) );
  DFFRX1 \key_reg[2]  ( .D(n328), .CK(n197), .RN(n132), .Q(key[2]) );
  DFFRX1 \key_reg[1]  ( .D(n329), .CK(n197), .RN(n132), .Q(key[1]) );
  DFFRX1 \key_reg[0]  ( .D(n330), .CK(n197), .RN(n132), .Q(key[0]) );
  DFFRX1 \din_reg[0]  ( .D(n274), .CK(n197), .RN(n132), .Q(din[0]) );
  DFFRX1 \din_reg[1]  ( .D(n273), .CK(n197), .RN(n131), .Q(din[1]) );
  DFFRX1 \din_reg[2]  ( .D(n272), .CK(n197), .RN(n131), .Q(din[2]) );
  DFFRX1 \din_reg[3]  ( .D(n271), .CK(n197), .RN(n131), .Q(din[3]) );
  DFFRX1 \din_reg[4]  ( .D(n270), .CK(n197), .RN(n131), .Q(din[4]) );
  DFFRX1 \din_reg[5]  ( .D(n269), .CK(n207), .RN(n131), .Q(din[5]) );
  DFFRX1 \din_reg[6]  ( .D(n268), .CK(n204), .RN(n131), .Q(din[6]) );
  DFFRX1 \din_reg[7]  ( .D(n267), .CK(n209), .RN(n131), .Q(din[7]) );
  DFFRX1 \din_reg[8]  ( .D(n266), .CK(n205), .RN(n131), .Q(din[8]) );
  DFFRX1 \din_reg[9]  ( .D(n265), .CK(n206), .RN(n131), .Q(din[9]) );
  DFFRX1 \din_reg[10]  ( .D(n264), .CK(n204), .RN(n130), .Q(din[10]) );
  DFFRX1 \din_reg[11]  ( .D(n263), .CK(n207), .RN(n130), .Q(din[11]) );
  DFFRX1 \din_reg[12]  ( .D(n262), .CK(n204), .RN(n130), .Q(din[12]) );
  DFFRX1 \din_reg[13]  ( .D(n261), .CK(n204), .RN(n130), .Q(din[13]) );
  DFFRX1 \din_reg[14]  ( .D(n260), .CK(n210), .RN(n130), .Q(din[14]) );
  DFFRX1 \din_reg[15]  ( .D(n259), .CK(n207), .RN(n130), .Q(din[15]) );
  DFFRX1 \din_reg[16]  ( .D(n258), .CK(n204), .RN(n130), .Q(din[16]) );
  DFFRX1 \din_reg[17]  ( .D(n257), .CK(n209), .RN(n130), .Q(din[17]) );
  DFFRX1 \din_reg[18]  ( .D(n256), .CK(n210), .RN(n130), .Q(din[18]) );
  DFFRX1 \din_reg[19]  ( .D(n255), .CK(n210), .RN(n129), .Q(din[19]) );
  DFFRX1 \din_reg[20]  ( .D(n254), .CK(n209), .RN(n129), .Q(din[20]) );
  DFFRX1 \din_reg[21]  ( .D(n253), .CK(n205), .RN(n129), .Q(din[21]) );
  DFFRX1 \din_reg[22]  ( .D(n252), .CK(n206), .RN(n129), .Q(din[22]) );
  DFFRX1 \din_reg[23]  ( .D(n251), .CK(n203), .RN(n129), .Q(din[23]) );
  DFFRX1 \din_reg[24]  ( .D(n250), .CK(n209), .RN(n129), .Q(din[24]) );
  DFFRX1 \din_reg[25]  ( .D(n249), .CK(n207), .RN(n129), .Q(din[25]) );
  DFFRX1 \din_reg[26]  ( .D(n248), .CK(n205), .RN(n129), .Q(din[26]) );
  DFFRX1 \din_reg[27]  ( .D(n247), .CK(n204), .RN(n129), .Q(din[27]) );
  DFFRX1 \din_reg[28]  ( .D(n246), .CK(n205), .RN(n142), .Q(din[28]) );
  DFFRX1 \din_reg[29]  ( .D(n245), .CK(n210), .RN(n143), .Q(din[29]) );
  DFFRX1 \din_reg[30]  ( .D(n244), .CK(n209), .RN(n144), .Q(din[30]) );
  DFFRX1 \din_reg[31]  ( .D(n243), .CK(n206), .RN(n145), .Q(din[31]) );
  DFFRX1 \din_reg[32]  ( .D(n242), .CK(n205), .RN(n144), .Q(din[32]) );
  DFFRX1 \din_reg[33]  ( .D(n241), .CK(n206), .RN(n139), .Q(din[33]) );
  DFFRX1 \din_reg[34]  ( .D(n240), .CK(n206), .RN(n140), .Q(din[34]) );
  DFFRX1 \din_reg[35]  ( .D(n239), .CK(n196), .RN(n142), .Q(din[35]) );
  DFFRX1 \din_reg[36]  ( .D(n238), .CK(n196), .RN(n145), .Q(din[36]) );
  DFFRX1 \din_reg[37]  ( .D(n237), .CK(n196), .RN(n145), .Q(din[37]) );
  DFFRX1 \din_reg[38]  ( .D(n236), .CK(n196), .RN(n143), .Q(din[38]) );
  DFFRX1 \din_reg[39]  ( .D(n235), .CK(n196), .RN(n144), .Q(din[39]) );
  DFFRX1 \din_reg[40]  ( .D(n234), .CK(n196), .RN(n139), .Q(din[40]) );
  DFFRX1 \din_reg[41]  ( .D(n233), .CK(n196), .RN(n145), .Q(din[41]) );
  DFFRX1 \din_reg[42]  ( .D(n232), .CK(n196), .RN(n139), .Q(din[42]) );
  DFFRX1 \din_reg[43]  ( .D(n231), .CK(n196), .RN(n140), .Q(din[43]) );
  DFFRX1 \din_reg[44]  ( .D(n230), .CK(n196), .RN(n141), .Q(din[44]) );
  DFFRX1 \din_reg[45]  ( .D(n229), .CK(n195), .RN(n144), .Q(din[45]) );
  DFFRX1 \din_reg[46]  ( .D(n228), .CK(n195), .RN(n128), .Q(din[46]) );
  DFFRX1 \din_reg[47]  ( .D(n227), .CK(n195), .RN(n145), .Q(din[47]) );
  DFFRX1 \din_reg[48]  ( .D(n226), .CK(n195), .RN(n140), .Q(din[48]) );
  DFFRX1 \din_reg[49]  ( .D(n225), .CK(n195), .RN(n139), .Q(din[49]) );
  DFFRX1 \din_reg[50]  ( .D(n224), .CK(n195), .RN(n140), .Q(din[50]) );
  DFFRX1 \din_reg[51]  ( .D(n223), .CK(n195), .RN(n141), .Q(din[51]) );
  DFFRX1 \din_reg[52]  ( .D(n222), .CK(n195), .RN(n142), .Q(din[52]) );
  DFFRX1 \din_reg[53]  ( .D(n221), .CK(n195), .RN(n143), .Q(din[53]) );
  DFFRX1 \din_reg[54]  ( .D(n220), .CK(n195), .RN(n143), .Q(din[54]) );
  DFFRX1 \din_reg[55]  ( .D(n219), .CK(clk), .RN(n140), .Q(din[55]) );
  DFFRX1 \din_reg[56]  ( .D(n218), .CK(clk), .RN(n141), .Q(din[56]) );
  DFFRX1 \din_reg[57]  ( .D(n217), .CK(clk), .RN(n142), .Q(din[57]) );
  DFFRX1 \din_reg[58]  ( .D(n216), .CK(clk), .RN(n143), .Q(din[58]) );
  DFFRX1 \din_reg[59]  ( .D(n215), .CK(clk), .RN(n145), .Q(din[59]) );
  DFFRX1 \din_reg[60]  ( .D(n214), .CK(n209), .RN(n144), .Q(din[60]) );
  DFFRX1 \din_reg[61]  ( .D(n213), .CK(n209), .RN(n128), .Q(din[61]) );
  DFFRX1 \din_reg[62]  ( .D(n212), .CK(n207), .RN(n141), .Q(din[62]) );
  DFFRX1 \din_reg[63]  ( .D(n211), .CK(clk), .RN(n128), .Q(din[63]) );
  DFFRX1 \cnt_reg[0]  ( .D(N10), .CK(n203), .RN(n138), .Q(cnt[0]) );
  DFFRX1 \cnt_reg[2]  ( .D(N12), .CK(n203), .RN(n138), .Q(cnt[2]) );
  DFFRX1 \cnt_reg[3]  ( .D(N13), .CK(n203), .RN(n138), .Q(cnt[3]) );
  CLKBUFX4 U3 ( .A(n176), .Y(n163) );
  CLKBUFX4 U4 ( .A(n176), .Y(n164) );
  AND2X2 U5 ( .A(reset_n), .B(desEnable), .Y(n128) );
  BUFX4 U6 ( .A(n143), .Y(n129) );
  BUFX4 U7 ( .A(n143), .Y(n130) );
  BUFX4 U8 ( .A(n142), .Y(n131) );
  BUFX4 U9 ( .A(n142), .Y(n132) );
  BUFX4 U10 ( .A(n141), .Y(n133) );
  BUFX4 U11 ( .A(n141), .Y(n134) );
  BUFX4 U12 ( .A(n140), .Y(n135) );
  BUFX4 U13 ( .A(n140), .Y(n136) );
  BUFX4 U14 ( .A(n210), .Y(n197) );
  BUFX4 U15 ( .A(n206), .Y(n198) );
  BUFX4 U16 ( .A(n206), .Y(n199) );
  BUFX4 U17 ( .A(n205), .Y(n200) );
  BUFX4 U18 ( .A(n205), .Y(n201) );
  BUFX4 U19 ( .A(n139), .Y(n137) );
  BUFX4 U20 ( .A(n139), .Y(n138) );
  BUFX4 U21 ( .A(n207), .Y(n195) );
  BUFX4 U22 ( .A(n207), .Y(n196) );
  BUFX4 U23 ( .A(n204), .Y(n202) );
  AOI222XL U24 ( .A0(desIn[62]), .A1(n188), .B0(n178), .B1(din[62]), .C0(
        desOut[62]), .C1(n154), .Y(n7) );
  AOI222XL U25 ( .A0(desIn[61]), .A1(n188), .B0(n168), .B1(din[61]), .C0(
        desOut[61]), .C1(n154), .Y(n8) );
  AOI222XL U26 ( .A0(desIn[60]), .A1(n188), .B0(n163), .B1(din[60]), .C0(
        desOut[60]), .C1(n154), .Y(n9) );
  AOI222XL U27 ( .A0(desIn[59]), .A1(n188), .B0(n176), .B1(din[59]), .C0(
        desOut[59]), .C1(n154), .Y(n10) );
  AOI222XL U28 ( .A0(desIn[58]), .A1(n188), .B0(n178), .B1(din[58]), .C0(
        desOut[58]), .C1(n154), .Y(n11) );
  AOI222XL U29 ( .A0(desIn[57]), .A1(n188), .B0(n177), .B1(din[57]), .C0(
        desOut[57]), .C1(n154), .Y(n12) );
  AOI222XL U30 ( .A0(desIn[56]), .A1(n188), .B0(n177), .B1(din[56]), .C0(
        desOut[56]), .C1(n154), .Y(n13) );
  AOI222XL U31 ( .A0(desIn[55]), .A1(n188), .B0(n174), .B1(din[55]), .C0(
        desOut[55]), .C1(n154), .Y(n14) );
  AOI222XL U32 ( .A0(desIn[54]), .A1(n187), .B0(n175), .B1(din[54]), .C0(
        desOut[54]), .C1(n154), .Y(n15) );
  AOI222XL U33 ( .A0(desIn[53]), .A1(n187), .B0(n178), .B1(din[53]), .C0(
        desOut[53]), .C1(n154), .Y(n16) );
  AOI222XL U34 ( .A0(desIn[52]), .A1(n187), .B0(n176), .B1(din[52]), .C0(
        desOut[52]), .C1(n153), .Y(n17) );
  AOI222XL U35 ( .A0(desIn[51]), .A1(n187), .B0(n172), .B1(din[51]), .C0(
        desOut[51]), .C1(n153), .Y(n18) );
  AOI222XL U36 ( .A0(desIn[50]), .A1(n187), .B0(n175), .B1(din[50]), .C0(
        desOut[50]), .C1(n153), .Y(n19) );
  AOI222XL U37 ( .A0(desIn[49]), .A1(n187), .B0(n173), .B1(din[49]), .C0(
        desOut[49]), .C1(n153), .Y(n20) );
  AOI222XL U38 ( .A0(desIn[48]), .A1(n187), .B0(n174), .B1(din[48]), .C0(
        desOut[48]), .C1(n153), .Y(n21) );
  AOI222XL U39 ( .A0(desIn[47]), .A1(n187), .B0(n173), .B1(din[47]), .C0(
        desOut[47]), .C1(n153), .Y(n22) );
  AOI222XL U40 ( .A0(desIn[46]), .A1(n187), .B0(n175), .B1(din[46]), .C0(
        desOut[46]), .C1(n153), .Y(n23) );
  AOI222XL U41 ( .A0(desIn[45]), .A1(n187), .B0(n173), .B1(din[45]), .C0(
        desOut[45]), .C1(n153), .Y(n24) );
  AOI222XL U42 ( .A0(desIn[44]), .A1(n186), .B0(n173), .B1(din[44]), .C0(
        desOut[44]), .C1(n153), .Y(n25) );
  AOI222XL U43 ( .A0(desIn[43]), .A1(n186), .B0(n178), .B1(din[43]), .C0(
        desOut[43]), .C1(n153), .Y(n26) );
  AOI222XL U44 ( .A0(desIn[42]), .A1(n186), .B0(n177), .B1(din[42]), .C0(
        desOut[42]), .C1(n152), .Y(n27) );
  AOI222XL U45 ( .A0(desIn[41]), .A1(n186), .B0(n164), .B1(din[41]), .C0(
        desOut[41]), .C1(n152), .Y(n28) );
  AOI222XL U46 ( .A0(desIn[40]), .A1(n186), .B0(n171), .B1(din[40]), .C0(
        desOut[40]), .C1(n152), .Y(n29) );
  AOI222XL U47 ( .A0(desIn[39]), .A1(n186), .B0(n163), .B1(din[39]), .C0(
        desOut[39]), .C1(n152), .Y(n30) );
  AOI222XL U48 ( .A0(desIn[38]), .A1(n186), .B0(n163), .B1(din[38]), .C0(
        desOut[38]), .C1(n152), .Y(n31) );
  AOI222XL U49 ( .A0(desIn[37]), .A1(n186), .B0(n163), .B1(din[37]), .C0(
        desOut[37]), .C1(n152), .Y(n32) );
  AOI222XL U50 ( .A0(desIn[36]), .A1(n186), .B0(n163), .B1(din[36]), .C0(
        desOut[36]), .C1(n152), .Y(n33) );
  AOI222XL U51 ( .A0(desIn[35]), .A1(n186), .B0(n163), .B1(din[35]), .C0(
        desOut[35]), .C1(n152), .Y(n34) );
  AOI222XL U52 ( .A0(desIn[34]), .A1(n185), .B0(n163), .B1(din[34]), .C0(
        desOut[34]), .C1(n152), .Y(n35) );
  AOI222XL U53 ( .A0(desIn[33]), .A1(n185), .B0(n163), .B1(din[33]), .C0(
        desOut[33]), .C1(n152), .Y(n36) );
  AOI222XL U54 ( .A0(desIn[32]), .A1(n185), .B0(n163), .B1(din[32]), .C0(
        desOut[32]), .C1(n151), .Y(n37) );
  AOI222XL U55 ( .A0(desIn[31]), .A1(n185), .B0(n164), .B1(din[31]), .C0(
        desOut[31]), .C1(n151), .Y(n38) );
  AOI222XL U56 ( .A0(desIn[30]), .A1(n185), .B0(n164), .B1(din[30]), .C0(
        desOut[30]), .C1(n151), .Y(n39) );
  AOI222XL U57 ( .A0(desIn[29]), .A1(n185), .B0(n164), .B1(din[29]), .C0(
        desOut[29]), .C1(n151), .Y(n40) );
  AOI222XL U58 ( .A0(desIn[28]), .A1(n185), .B0(n164), .B1(din[28]), .C0(
        desOut[28]), .C1(n151), .Y(n41) );
  AOI222XL U59 ( .A0(desIn[27]), .A1(n185), .B0(n164), .B1(din[27]), .C0(
        desOut[27]), .C1(n151), .Y(n42) );
  AOI222XL U60 ( .A0(desIn[26]), .A1(n185), .B0(n164), .B1(din[26]), .C0(
        desOut[26]), .C1(n151), .Y(n43) );
  AOI222XL U61 ( .A0(desIn[25]), .A1(n185), .B0(n164), .B1(din[25]), .C0(
        desOut[25]), .C1(n151), .Y(n44) );
  AOI222XL U62 ( .A0(desIn[24]), .A1(n184), .B0(n164), .B1(din[24]), .C0(
        desOut[24]), .C1(n151), .Y(n45) );
  AOI222XL U63 ( .A0(desIn[23]), .A1(n184), .B0(n165), .B1(din[23]), .C0(
        desOut[23]), .C1(n151), .Y(n46) );
  AOI222XL U64 ( .A0(desIn[22]), .A1(n184), .B0(n165), .B1(din[22]), .C0(
        desOut[22]), .C1(n150), .Y(n47) );
  AOI222XL U65 ( .A0(desIn[21]), .A1(n184), .B0(n165), .B1(din[21]), .C0(
        desOut[21]), .C1(n150), .Y(n48) );
  AOI222XL U66 ( .A0(desIn[20]), .A1(n184), .B0(n165), .B1(din[20]), .C0(
        desOut[20]), .C1(n150), .Y(n49) );
  AOI222XL U67 ( .A0(desIn[19]), .A1(n184), .B0(n165), .B1(din[19]), .C0(
        desOut[19]), .C1(n150), .Y(n50) );
  AOI222XL U68 ( .A0(desIn[18]), .A1(n184), .B0(n165), .B1(din[18]), .C0(
        desOut[18]), .C1(n150), .Y(n51) );
  AOI222XL U69 ( .A0(desIn[17]), .A1(n184), .B0(n165), .B1(din[17]), .C0(
        desOut[17]), .C1(n150), .Y(n52) );
  AOI222XL U70 ( .A0(desIn[16]), .A1(n184), .B0(n165), .B1(din[16]), .C0(
        desOut[16]), .C1(n150), .Y(n53) );
  AOI222XL U71 ( .A0(desIn[15]), .A1(n184), .B0(n166), .B1(din[15]), .C0(
        desOut[15]), .C1(n150), .Y(n54) );
  AOI222XL U72 ( .A0(desIn[14]), .A1(n183), .B0(n166), .B1(din[14]), .C0(
        desOut[14]), .C1(n150), .Y(n55) );
  AOI222XL U73 ( .A0(desIn[13]), .A1(n183), .B0(n166), .B1(din[13]), .C0(
        desOut[13]), .C1(n150), .Y(n56) );
  AOI222XL U74 ( .A0(desIn[12]), .A1(n183), .B0(n166), .B1(din[12]), .C0(
        desOut[12]), .C1(n149), .Y(n57) );
  AOI222XL U75 ( .A0(desIn[11]), .A1(n183), .B0(n166), .B1(din[11]), .C0(
        desOut[11]), .C1(n149), .Y(n58) );
  AOI222XL U76 ( .A0(desIn[10]), .A1(n183), .B0(n166), .B1(din[10]), .C0(
        desOut[10]), .C1(n149), .Y(n59) );
  AOI222XL U77 ( .A0(desIn[9]), .A1(n183), .B0(n166), .B1(din[9]), .C0(
        desOut[9]), .C1(n149), .Y(n60) );
  AOI222XL U78 ( .A0(desIn[8]), .A1(n183), .B0(n166), .B1(din[8]), .C0(
        desOut[8]), .C1(n149), .Y(n61) );
  AOI222XL U79 ( .A0(desIn[7]), .A1(n183), .B0(n167), .B1(din[7]), .C0(
        desOut[7]), .C1(n149), .Y(n62) );
  AOI222XL U80 ( .A0(desIn[6]), .A1(n183), .B0(n167), .B1(din[6]), .C0(
        desOut[6]), .C1(n149), .Y(n63) );
  AOI222XL U81 ( .A0(desIn[5]), .A1(n183), .B0(n167), .B1(din[5]), .C0(
        desOut[5]), .C1(n149), .Y(n64) );
  AOI222XL U82 ( .A0(desIn[4]), .A1(n182), .B0(n167), .B1(din[4]), .C0(
        desOut[4]), .C1(n149), .Y(n65) );
  AOI222XL U83 ( .A0(desIn[3]), .A1(n182), .B0(n167), .B1(din[3]), .C0(
        desOut[3]), .C1(n149), .Y(n66) );
  AOI222XL U84 ( .A0(desIn[2]), .A1(n182), .B0(n167), .B1(din[2]), .C0(
        desOut[2]), .C1(n148), .Y(n67) );
  AOI222XL U85 ( .A0(desIn[1]), .A1(n182), .B0(n167), .B1(din[1]), .C0(
        desOut[1]), .C1(n148), .Y(n68) );
  AOI222XL U86 ( .A0(desIn[0]), .A1(n182), .B0(n167), .B1(din[0]), .C0(
        desOut[0]), .C1(n148), .Y(n69) );
  AOI222XL U87 ( .A0(key1[44]), .A1(n181), .B0(n169), .B1(key[44]), .C0(
        key2[44]), .C1(n147), .Y(n81) );
  AOI222XL U88 ( .A0(key1[45]), .A1(n181), .B0(n169), .B1(key[45]), .C0(
        key2[45]), .C1(n147), .Y(n80) );
  AOI222XL U89 ( .A0(key1[46]), .A1(n181), .B0(n169), .B1(key[46]), .C0(
        key2[46]), .C1(n147), .Y(n79) );
  AOI222XL U90 ( .A0(key1[47]), .A1(n181), .B0(n169), .B1(key[47]), .C0(
        key2[47]), .C1(n147), .Y(n78) );
  AOI222XL U91 ( .A0(desIn[63]), .A1(n193), .B0(n176), .B1(din[63]), .C0(
        desOut[63]), .C1(n155), .Y(n4) );
  AOI222XL U92 ( .A0(key1[0]), .A1(n194), .B0(n165), .B1(key[0]), .C0(key2[0]), 
        .C1(n155), .Y(n125) );
  AOI222XL U93 ( .A0(key1[1]), .A1(n194), .B0(n175), .B1(key[1]), .C0(key2[1]), 
        .C1(n155), .Y(n124) );
  AOI222XL U94 ( .A0(key1[2]), .A1(n189), .B0(n173), .B1(key[2]), .C0(key2[2]), 
        .C1(n156), .Y(n123) );
  AOI222XL U95 ( .A0(key1[3]), .A1(n190), .B0(n166), .B1(key[3]), .C0(key2[3]), 
        .C1(n161), .Y(n122) );
  AOI222XL U96 ( .A0(key1[4]), .A1(n189), .B0(n178), .B1(key[4]), .C0(key2[4]), 
        .C1(n159), .Y(n121) );
  AOI222XL U97 ( .A0(key1[5]), .A1(n192), .B0(n177), .B1(key[5]), .C0(key2[5]), 
        .C1(n156), .Y(n120) );
  AOI222XL U98 ( .A0(key1[6]), .A1(n191), .B0(n163), .B1(key[6]), .C0(key2[6]), 
        .C1(n157), .Y(n119) );
  AOI222XL U99 ( .A0(key1[7]), .A1(n192), .B0(n174), .B1(key[7]), .C0(key2[7]), 
        .C1(n158), .Y(n118) );
  AOI222XL U100 ( .A0(key1[8]), .A1(N3), .B0(n170), .B1(key[8]), .C0(key2[8]), 
        .C1(n160), .Y(n117) );
  AOI222XL U101 ( .A0(key1[9]), .A1(n193), .B0(n174), .B1(key[9]), .C0(key2[9]), .C1(n157), .Y(n116) );
  AOI222XL U102 ( .A0(key1[10]), .A1(n191), .B0(n175), .B1(key[10]), .C0(
        key2[10]), .C1(n156), .Y(n115) );
  AOI222XL U103 ( .A0(key1[11]), .A1(n190), .B0(n177), .B1(key[11]), .C0(
        key2[11]), .C1(n157), .Y(n114) );
  AOI222XL U104 ( .A0(key1[12]), .A1(n193), .B0(n178), .B1(key[12]), .C0(
        key2[12]), .C1(n160), .Y(n113) );
  AOI222XL U105 ( .A0(key1[13]), .A1(n192), .B0(n169), .B1(key[13]), .C0(
        key2[13]), .C1(n156), .Y(n112) );
  AOI222XL U106 ( .A0(key1[14]), .A1(n189), .B0(n164), .B1(key[14]), .C0(
        key2[14]), .C1(n157), .Y(n111) );
  AOI222XL U107 ( .A0(key1[15]), .A1(n193), .B0(n174), .B1(key[15]), .C0(
        key2[15]), .C1(n158), .Y(n110) );
  AOI222XL U108 ( .A0(key1[16]), .A1(n194), .B0(n172), .B1(key[16]), .C0(
        key2[16]), .C1(n160), .Y(n109) );
  AOI222XL U109 ( .A0(key1[17]), .A1(N3), .B0(n172), .B1(key[17]), .C0(
        key2[17]), .C1(n159), .Y(n108) );
  AOI222XL U110 ( .A0(key1[18]), .A1(n190), .B0(n172), .B1(key[18]), .C0(
        key2[18]), .C1(n162), .Y(n107) );
  AOI222XL U111 ( .A0(key1[19]), .A1(n191), .B0(n172), .B1(key[19]), .C0(
        key2[19]), .C1(n159), .Y(n106) );
  AOI222XL U112 ( .A0(key1[20]), .A1(n179), .B0(n172), .B1(key[20]), .C0(
        key2[20]), .C1(n162), .Y(n105) );
  AOI222XL U113 ( .A0(key1[21]), .A1(n194), .B0(n172), .B1(key[21]), .C0(
        key2[21]), .C1(n162), .Y(n104) );
  AOI222XL U114 ( .A0(key1[22]), .A1(n179), .B0(n172), .B1(key[22]), .C0(
        key2[22]), .C1(n155), .Y(n103) );
  AOI222XL U115 ( .A0(key1[23]), .A1(n179), .B0(n172), .B1(key[23]), .C0(
        key2[23]), .C1(n162), .Y(n102) );
  AOI222XL U116 ( .A0(key1[24]), .A1(n179), .B0(n171), .B1(key[24]), .C0(
        key2[24]), .C1(n162), .Y(n101) );
  AOI222XL U117 ( .A0(key1[25]), .A1(n182), .B0(n171), .B1(key[25]), .C0(
        key2[25]), .C1(n155), .Y(n100) );
  AOI222XL U118 ( .A0(key1[26]), .A1(n179), .B0(n171), .B1(key[26]), .C0(
        key2[26]), .C1(n158), .Y(n99) );
  AOI222XL U119 ( .A0(key1[27]), .A1(n179), .B0(n171), .B1(key[27]), .C0(
        key2[27]), .C1(n161), .Y(n98) );
  AOI222XL U120 ( .A0(key1[28]), .A1(n179), .B0(n171), .B1(key[28]), .C0(
        key2[28]), .C1(n162), .Y(n97) );
  AOI222XL U121 ( .A0(key1[29]), .A1(n179), .B0(n171), .B1(key[29]), .C0(
        key2[29]), .C1(n146), .Y(n96) );
  AOI222XL U122 ( .A0(key1[30]), .A1(n179), .B0(n171), .B1(key[30]), .C0(
        key2[30]), .C1(n146), .Y(n95) );
  AOI222XL U123 ( .A0(key1[31]), .A1(n179), .B0(n171), .B1(key[31]), .C0(
        key2[31]), .C1(n146), .Y(n94) );
  AOI222XL U124 ( .A0(key1[32]), .A1(n180), .B0(n170), .B1(key[32]), .C0(
        key2[32]), .C1(n146), .Y(n93) );
  AOI222XL U125 ( .A0(key1[33]), .A1(n180), .B0(n170), .B1(key[33]), .C0(
        key2[33]), .C1(n146), .Y(n92) );
  AOI222XL U126 ( .A0(key1[34]), .A1(n180), .B0(n170), .B1(key[34]), .C0(
        key2[34]), .C1(n146), .Y(n91) );
  AOI222XL U127 ( .A0(key1[35]), .A1(n180), .B0(n170), .B1(key[35]), .C0(
        key2[35]), .C1(n146), .Y(n90) );
  AOI222XL U128 ( .A0(key1[36]), .A1(n180), .B0(n170), .B1(key[36]), .C0(
        key2[36]), .C1(n146), .Y(n89) );
  AOI222XL U129 ( .A0(key1[37]), .A1(n180), .B0(n170), .B1(key[37]), .C0(
        key2[37]), .C1(n146), .Y(n88) );
  AOI222XL U130 ( .A0(key1[38]), .A1(n180), .B0(n170), .B1(key[38]), .C0(
        key2[38]), .C1(n146), .Y(n87) );
  AOI222XL U131 ( .A0(key1[39]), .A1(n180), .B0(n170), .B1(key[39]), .C0(
        key2[39]), .C1(n147), .Y(n86) );
  AOI222XL U132 ( .A0(key1[40]), .A1(n180), .B0(n169), .B1(key[40]), .C0(
        key2[40]), .C1(n147), .Y(n85) );
  AOI222XL U133 ( .A0(key1[41]), .A1(n180), .B0(n169), .B1(key[41]), .C0(
        key2[41]), .C1(n147), .Y(n84) );
  AOI222XL U134 ( .A0(key1[42]), .A1(n181), .B0(n169), .B1(key[42]), .C0(
        key2[42]), .C1(n147), .Y(n83) );
  AOI222XL U135 ( .A0(key1[43]), .A1(n181), .B0(n169), .B1(key[43]), .C0(
        key2[43]), .C1(n147), .Y(n82) );
  AOI222XL U136 ( .A0(key1[48]), .A1(n181), .B0(n168), .B1(key[48]), .C0(
        key2[48]), .C1(n147), .Y(n77) );
  AOI222XL U137 ( .A0(key1[49]), .A1(n181), .B0(n168), .B1(key[49]), .C0(
        key2[49]), .C1(n148), .Y(n76) );
  AOI222XL U138 ( .A0(key1[50]), .A1(n181), .B0(n168), .B1(key[50]), .C0(
        key2[50]), .C1(n148), .Y(n75) );
  AOI222XL U139 ( .A0(key1[51]), .A1(n181), .B0(n168), .B1(key[51]), .C0(
        key2[51]), .C1(n148), .Y(n74) );
  AOI222XL U140 ( .A0(key1[52]), .A1(n182), .B0(n168), .B1(key[52]), .C0(
        key2[52]), .C1(n148), .Y(n73) );
  AOI222XL U141 ( .A0(key1[53]), .A1(n182), .B0(n168), .B1(key[53]), .C0(
        key2[53]), .C1(n148), .Y(n72) );
  AOI222XL U142 ( .A0(key1[54]), .A1(n182), .B0(n168), .B1(key[54]), .C0(
        key2[54]), .C1(n148), .Y(n71) );
  AOI222XL U143 ( .A0(key1[55]), .A1(n182), .B0(n168), .B1(key[55]), .C0(
        key2[55]), .C1(n148), .Y(n70) );
  BUFX4 U144 ( .A(n5), .Y(n165) );
  BUFX4 U145 ( .A(n167), .Y(n166) );
  BUFX4 U146 ( .A(n175), .Y(n167) );
  BUFX4 U147 ( .A(n173), .Y(n172) );
  BUFX4 U148 ( .A(n173), .Y(n171) );
  BUFX4 U149 ( .A(n174), .Y(n170) );
  BUFX4 U150 ( .A(n174), .Y(n169) );
  BUFX4 U151 ( .A(n175), .Y(n168) );
  CLKBUFX3 U152 ( .A(n5), .Y(n176) );
  CLKBUFX3 U153 ( .A(n178), .Y(n173) );
  CLKBUFX3 U154 ( .A(n177), .Y(n174) );
  CLKBUFX3 U155 ( .A(n177), .Y(n175) );
  CLKBUFX3 U156 ( .A(n176), .Y(n178) );
  CLKBUFX3 U157 ( .A(n176), .Y(n177) );
  CLKBUFX6 U158 ( .A(n190), .Y(n186) );
  CLKBUFX6 U159 ( .A(n190), .Y(n185) );
  CLKBUFX6 U160 ( .A(n194), .Y(n184) );
  CLKBUFX6 U161 ( .A(n194), .Y(n183) );
  CLKBUFX6 U162 ( .A(n192), .Y(n179) );
  CLKBUFX6 U163 ( .A(n192), .Y(n180) );
  CLKBUFX6 U164 ( .A(n191), .Y(n181) );
  CLKBUFX6 U165 ( .A(n191), .Y(n182) );
  CLKBUFX6 U166 ( .A(n157), .Y(n153) );
  CLKBUFX6 U167 ( .A(n157), .Y(n152) );
  CLKBUFX6 U168 ( .A(n158), .Y(n151) );
  CLKBUFX6 U169 ( .A(n158), .Y(n150) );
  CLKBUFX6 U170 ( .A(n159), .Y(n149) );
  CLKBUFX6 U171 ( .A(n160), .Y(n146) );
  CLKBUFX6 U172 ( .A(n160), .Y(n147) );
  CLKBUFX6 U173 ( .A(n159), .Y(n148) );
  CLKBUFX6 U174 ( .A(n189), .Y(n187) );
  CLKBUFX6 U175 ( .A(n156), .Y(n154) );
  BUFX4 U176 ( .A(n189), .Y(n188) );
  CLKBUFX3 U177 ( .A(n155), .Y(n157) );
  CLKBUFX3 U178 ( .A(n191), .Y(n190) );
  CLKBUFX3 U179 ( .A(n6), .Y(n158) );
  CLKBUFX3 U180 ( .A(n193), .Y(n192) );
  CLKBUFX3 U181 ( .A(n161), .Y(n160) );
  CLKBUFX3 U182 ( .A(n193), .Y(n191) );
  CLKBUFX3 U183 ( .A(n161), .Y(n159) );
  NOR2X1 U184 ( .A(n161), .B(n189), .Y(n5) );
  CLKBUFX3 U185 ( .A(N3), .Y(n193) );
  CLKBUFX3 U186 ( .A(n6), .Y(n161) );
  CLKBUFX3 U187 ( .A(n141), .Y(n143) );
  CLKBUFX3 U188 ( .A(n139), .Y(n142) );
  CLKBUFX3 U189 ( .A(n144), .Y(n141) );
  CLKBUFX3 U190 ( .A(n144), .Y(n140) );
  CLKBUFX3 U191 ( .A(n208), .Y(n206) );
  CLKBUFX3 U192 ( .A(n208), .Y(n205) );
  CLKBUFX3 U193 ( .A(n162), .Y(n156) );
  CLKBUFX3 U194 ( .A(n158), .Y(n162) );
  CLKBUFX3 U195 ( .A(n194), .Y(n189) );
  CLKBUFX3 U196 ( .A(n192), .Y(n194) );
  CLKBUFX3 U197 ( .A(n204), .Y(n203) );
  NAND2BX1 U198 ( .AN(N7), .B(n193), .Y(N12) );
  CLKBUFX3 U199 ( .A(n128), .Y(n144) );
  AND2X2 U200 ( .A(N8), .B(n191), .Y(N13) );
  AND2X2 U201 ( .A(N6), .B(n190), .Y(N11) );
  CLKBUFX3 U202 ( .A(n210), .Y(n208) );
  CLKBUFX3 U203 ( .A(clk), .Y(n207) );
  CLKBUFX3 U204 ( .A(n145), .Y(n139) );
  CLKBUFX3 U205 ( .A(n128), .Y(n145) );
  CLKBUFX3 U206 ( .A(n209), .Y(n204) );
  CLKBUFX3 U207 ( .A(n210), .Y(n209) );
  NAND2X1 U208 ( .A(n126), .B(n190), .Y(n127) );
  AOI2BB1X1 U209 ( .A0N(cnt[3]), .A1N(cnt[2]), .B0(n2), .Y(n1) );
  CLKINVX1 U210 ( .A(n1), .Y(N3) );
  NAND2X1 U211 ( .A(n3), .B(n189), .Y(N14) );
  XNOR2X1 U212 ( .A(\add_24/carry[4] ), .B(cnt[4]), .Y(n3) );
  NAND2X1 U213 ( .A(cnt[0]), .B(n192), .Y(N10) );
  CLKBUFX3 U214 ( .A(clk), .Y(n210) );
  NOR2BX1 U215 ( .AN(n126), .B(N3), .Y(n6) );
  CLKINVX1 U216 ( .A(n4), .Y(n211) );
  CLKBUFX3 U217 ( .A(n156), .Y(n155) );
  CLKINVX1 U218 ( .A(n7), .Y(n212) );
  CLKINVX1 U219 ( .A(n8), .Y(n213) );
  CLKINVX1 U220 ( .A(n9), .Y(n214) );
  CLKINVX1 U221 ( .A(n10), .Y(n215) );
  CLKINVX1 U222 ( .A(n11), .Y(n216) );
  CLKINVX1 U223 ( .A(n12), .Y(n217) );
  CLKINVX1 U224 ( .A(n13), .Y(n218) );
  CLKINVX1 U225 ( .A(n14), .Y(n219) );
  CLKINVX1 U226 ( .A(n15), .Y(n220) );
  CLKINVX1 U227 ( .A(n16), .Y(n221) );
  CLKINVX1 U228 ( .A(n17), .Y(n222) );
  CLKINVX1 U229 ( .A(n18), .Y(n223) );
  CLKINVX1 U230 ( .A(n19), .Y(n224) );
  CLKINVX1 U231 ( .A(n20), .Y(n225) );
  CLKINVX1 U232 ( .A(n21), .Y(n226) );
  CLKINVX1 U233 ( .A(n22), .Y(n227) );
  CLKINVX1 U234 ( .A(n23), .Y(n228) );
  CLKINVX1 U235 ( .A(n24), .Y(n229) );
  CLKINVX1 U236 ( .A(n25), .Y(n230) );
  CLKINVX1 U237 ( .A(n26), .Y(n231) );
  CLKINVX1 U238 ( .A(n27), .Y(n232) );
  CLKINVX1 U239 ( .A(n28), .Y(n233) );
  CLKINVX1 U240 ( .A(n29), .Y(n234) );
  CLKINVX1 U241 ( .A(n30), .Y(n235) );
  CLKINVX1 U242 ( .A(n31), .Y(n236) );
  CLKINVX1 U243 ( .A(n32), .Y(n237) );
  CLKINVX1 U244 ( .A(n33), .Y(n238) );
  CLKINVX1 U245 ( .A(n34), .Y(n239) );
  CLKINVX1 U246 ( .A(n35), .Y(n240) );
  CLKINVX1 U247 ( .A(n36), .Y(n241) );
  CLKINVX1 U248 ( .A(n37), .Y(n242) );
  CLKINVX1 U249 ( .A(n38), .Y(n243) );
  CLKINVX1 U250 ( .A(n39), .Y(n244) );
  CLKINVX1 U251 ( .A(n40), .Y(n245) );
  CLKINVX1 U252 ( .A(n41), .Y(n246) );
  CLKINVX1 U253 ( .A(n42), .Y(n247) );
  CLKINVX1 U254 ( .A(n43), .Y(n248) );
  CLKINVX1 U255 ( .A(n44), .Y(n249) );
  CLKINVX1 U256 ( .A(n45), .Y(n250) );
  CLKINVX1 U257 ( .A(n46), .Y(n251) );
  CLKINVX1 U258 ( .A(n47), .Y(n252) );
  CLKINVX1 U259 ( .A(n48), .Y(n253) );
  CLKINVX1 U260 ( .A(n49), .Y(n254) );
  CLKINVX1 U261 ( .A(n50), .Y(n255) );
  CLKINVX1 U262 ( .A(n51), .Y(n256) );
  CLKINVX1 U263 ( .A(n52), .Y(n257) );
  CLKINVX1 U264 ( .A(n53), .Y(n258) );
  CLKINVX1 U265 ( .A(n54), .Y(n259) );
  CLKINVX1 U266 ( .A(n55), .Y(n260) );
  CLKINVX1 U267 ( .A(n56), .Y(n261) );
  CLKINVX1 U268 ( .A(n57), .Y(n262) );
  CLKINVX1 U269 ( .A(n58), .Y(n263) );
  CLKINVX1 U270 ( .A(n59), .Y(n264) );
  CLKINVX1 U271 ( .A(n60), .Y(n265) );
  CLKINVX1 U272 ( .A(n61), .Y(n266) );
  CLKINVX1 U273 ( .A(n62), .Y(n267) );
  CLKINVX1 U274 ( .A(n63), .Y(n268) );
  CLKINVX1 U275 ( .A(n64), .Y(n269) );
  CLKINVX1 U276 ( .A(n65), .Y(n270) );
  CLKINVX1 U277 ( .A(n66), .Y(n271) );
  CLKINVX1 U278 ( .A(n67), .Y(n272) );
  CLKINVX1 U279 ( .A(n68), .Y(n273) );
  CLKINVX1 U280 ( .A(n69), .Y(n274) );
  CLKINVX1 U281 ( .A(n81), .Y(n286) );
  CLKINVX1 U282 ( .A(n80), .Y(n285) );
  CLKINVX1 U283 ( .A(n79), .Y(n284) );
  CLKINVX1 U284 ( .A(n78), .Y(n283) );
  CLKINVX1 U285 ( .A(n125), .Y(n330) );
  CLKINVX1 U286 ( .A(n124), .Y(n329) );
  CLKINVX1 U287 ( .A(n123), .Y(n328) );
  CLKINVX1 U288 ( .A(n122), .Y(n327) );
  CLKINVX1 U289 ( .A(n121), .Y(n326) );
  CLKINVX1 U290 ( .A(n120), .Y(n325) );
  CLKINVX1 U291 ( .A(n119), .Y(n324) );
  CLKINVX1 U292 ( .A(n118), .Y(n323) );
  CLKINVX1 U293 ( .A(n117), .Y(n322) );
  CLKINVX1 U294 ( .A(n116), .Y(n321) );
  CLKINVX1 U295 ( .A(n115), .Y(n320) );
  CLKINVX1 U296 ( .A(n114), .Y(n319) );
  CLKINVX1 U297 ( .A(n113), .Y(n318) );
  CLKINVX1 U298 ( .A(n112), .Y(n317) );
  CLKINVX1 U299 ( .A(n111), .Y(n316) );
  CLKINVX1 U300 ( .A(n110), .Y(n315) );
  CLKINVX1 U301 ( .A(n109), .Y(n314) );
  CLKINVX1 U302 ( .A(n108), .Y(n313) );
  CLKINVX1 U303 ( .A(n107), .Y(n312) );
  CLKINVX1 U304 ( .A(n106), .Y(n311) );
  CLKINVX1 U305 ( .A(n105), .Y(n310) );
  CLKINVX1 U306 ( .A(n104), .Y(n309) );
  CLKINVX1 U307 ( .A(n103), .Y(n308) );
  CLKINVX1 U308 ( .A(n102), .Y(n307) );
  CLKINVX1 U309 ( .A(n101), .Y(n306) );
  CLKINVX1 U310 ( .A(n100), .Y(n305) );
  CLKINVX1 U311 ( .A(n99), .Y(n304) );
  CLKINVX1 U312 ( .A(n98), .Y(n303) );
  CLKINVX1 U313 ( .A(n97), .Y(n302) );
  CLKINVX1 U314 ( .A(n96), .Y(n301) );
  CLKINVX1 U315 ( .A(n95), .Y(n300) );
  CLKINVX1 U316 ( .A(n94), .Y(n299) );
  CLKINVX1 U317 ( .A(n93), .Y(n298) );
  CLKINVX1 U318 ( .A(n92), .Y(n297) );
  CLKINVX1 U319 ( .A(n91), .Y(n296) );
  CLKINVX1 U320 ( .A(n90), .Y(n295) );
  CLKINVX1 U321 ( .A(n89), .Y(n294) );
  CLKINVX1 U322 ( .A(n88), .Y(n293) );
  CLKINVX1 U323 ( .A(n87), .Y(n292) );
  CLKINVX1 U324 ( .A(n86), .Y(n291) );
  CLKINVX1 U325 ( .A(n85), .Y(n290) );
  CLKINVX1 U326 ( .A(n84), .Y(n289) );
  CLKINVX1 U327 ( .A(n83), .Y(n288) );
  CLKINVX1 U328 ( .A(n82), .Y(n287) );
  CLKINVX1 U329 ( .A(n77), .Y(n282) );
  CLKINVX1 U330 ( .A(n76), .Y(n281) );
  CLKINVX1 U331 ( .A(n75), .Y(n280) );
  CLKINVX1 U332 ( .A(n74), .Y(n279) );
  CLKINVX1 U333 ( .A(n73), .Y(n278) );
  CLKINVX1 U334 ( .A(n72), .Y(n277) );
  CLKINVX1 U335 ( .A(n71), .Y(n276) );
  CLKINVX1 U336 ( .A(n70), .Y(n275) );
endmodule


module seg_decoder_DW01_inc_0 ( A, SUM );
  input [12:0] A;
  output [12:0] SUM;

  wire   [12:2] carry;

  ADDHXL U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXL U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDHXL U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHXL U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  XOR2X1 U1 ( .A(carry[12]), .B(A[12]), .Y(SUM[12]) );
  CLKINVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module seg_decoder ( desOut, desEnable, reset_n, clk, segout1, segout2 );
  input [64:1] desOut;
  output [6:0] segout1;
  output [6:0] segout2;
  input desEnable, reset_n, clk;
  wire   N240, N241, N242, N243, N244, N245, N246, N247, N248, N249, N250,
         N251, N252, n7, n8, n10, n12, n14, n16, n17, n18, n21, n22, n23, n25,
         n26, n28, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n1, n2, n3, n4, n5, n6, n9,
         n11, n13, n15, n19, n20, n24, n27, n29, n53, n151, n152, n153, n154,
         n155, n156, n157;
  wire   [3:0] i_hex;
  wire   [4:0] decoderin1;
  wire   [4:0] decoderin2;
  wire   [13:1] clk_div;
  wire   [1:0] i_idle;
  wire   [1:0] state;

  DFFRX4 \i_hex_reg[0]  ( .D(n149), .CK(n5), .RN(n157), .Q(i_hex[0]), .QN(n23)
         );
  DFFRX4 \i_hex_reg[3]  ( .D(n148), .CK(n5), .RN(n157), .Q(i_hex[3]), .QN(n18)
         );
  DFFRX4 \i_hex_reg[1]  ( .D(n143), .CK(n5), .RN(n157), .Q(i_hex[1]), .QN(n22)
         );
  DFFRX4 \i_hex_reg[2]  ( .D(n142), .CK(n5), .RN(n157), .Q(i_hex[2]), .QN(n21)
         );
  DFFRX4 \decoderin2_reg[3]  ( .D(decoderin1[3]), .CK(n5), .RN(n157), .Q(
        decoderin2[3]), .QN(n26) );
  DFFRX4 \decoderin2_reg[2]  ( .D(decoderin1[2]), .CK(n5), .RN(n157), .Q(
        decoderin2[2]), .QN(n28) );
  DFFRX4 \decoderin2_reg[1]  ( .D(decoderin1[1]), .CK(n5), .RN(n157), .Q(
        decoderin2[1]), .QN(n30) );
  NOR4X2 U23 ( .A(n25), .B(decoderin2[1]), .C(decoderin2[2]), .D(decoderin2[3]), .Y(n39) );
  NOR2X2 U24 ( .A(n31), .B(decoderin2[3]), .Y(n35) );
  NAND2X2 U27 ( .A(decoderin2[1]), .B(n28), .Y(n37) );
  NAND2X2 U28 ( .A(decoderin2[2]), .B(n30), .Y(n36) );
  NOR2X2 U52 ( .A(n17), .B(decoderin1[3]), .Y(n55) );
  NOR2X2 U55 ( .A(n54), .B(decoderin1[0]), .Y(n61) );
  NAND2X2 U56 ( .A(decoderin1[2]), .B(n16), .Y(n54) );
  NOR3BX2 U93 ( .AN(n121), .B(n21), .C(n22), .Y(n80) );
  NOR3BX2 U95 ( .AN(n122), .B(n18), .C(n23), .Y(n77) );
  NOR3X2 U98 ( .A(n18), .B(n22), .C(n124), .Y(n85) );
  NOR3BX2 U99 ( .AN(n121), .B(n22), .C(i_hex[2]), .Y(n84) );
  NOR3BX2 U100 ( .AN(n121), .B(i_hex[1]), .C(i_hex[2]), .Y(n82) );
  NOR2X2 U101 ( .A(n18), .B(i_hex[0]), .Y(n121) );
  NOR3BX2 U105 ( .AN(n127), .B(n21), .C(i_hex[0]), .Y(n89) );
  NOR3BX2 U106 ( .AN(n122), .B(i_hex[0]), .C(i_hex[3]), .Y(n87) );
  NOR3BX2 U107 ( .AN(n122), .B(n23), .C(i_hex[3]), .Y(n86) );
  NOR2X2 U108 ( .A(n21), .B(i_hex[1]), .Y(n122) );
  NOR2BX2 U111 ( .AN(n127), .B(n124), .Y(n94) );
  NOR3BX2 U112 ( .AN(n127), .B(i_hex[0]), .C(i_hex[2]), .Y(n93) );
  NOR3X2 U114 ( .A(i_hex[1]), .B(i_hex[3]), .C(n124), .Y(n90) );
  NAND2X2 U115 ( .A(state[1]), .B(state[0]), .Y(n71) );
  NOR2X2 U133 ( .A(n22), .B(i_hex[3]), .Y(n127) );
  NAND2X2 U135 ( .A(state[0]), .B(n7), .Y(n129) );
  DFFSX4 \decoderin2_reg[4]  ( .D(decoderin1[4]), .CK(n4), .SN(n2), .Q(
        decoderin2[4]), .QN(n25) );
  DFFSX4 \decoderin2_reg[0]  ( .D(decoderin1[0]), .CK(n5), .SN(n157), .Q(
        decoderin2[0]), .QN(n31) );
  seg_decoder_DW01_inc_0 add_124 ( .A({n4, clk_div[12:1]}), .SUM({N252, N251, 
        N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240}) );
  DFFRX2 \state_reg[1]  ( .D(n147), .CK(n4), .RN(n2), .Q(state[1]), .QN(n7) );
  DFFRX1 \clk_div_reg[2]  ( .D(N241), .CK(n9), .RN(reset_n), .Q(clk_div[2]) );
  DFFRX1 \clk_div_reg[3]  ( .D(N242), .CK(n9), .RN(reset_n), .Q(clk_div[3]) );
  DFFRX1 \clk_div_reg[4]  ( .D(N243), .CK(n9), .RN(n11), .Q(clk_div[4]) );
  DFFRX1 \clk_div_reg[5]  ( .D(N244), .CK(n6), .RN(n11), .Q(clk_div[5]) );
  DFFRX1 \clk_div_reg[6]  ( .D(N245), .CK(n6), .RN(n11), .Q(clk_div[6]) );
  DFFRX1 \clk_div_reg[7]  ( .D(N246), .CK(n6), .RN(n11), .Q(clk_div[7]) );
  DFFRX1 \clk_div_reg[8]  ( .D(N247), .CK(n6), .RN(n11), .Q(clk_div[8]) );
  DFFRX1 \clk_div_reg[9]  ( .D(N248), .CK(n6), .RN(n11), .Q(clk_div[9]) );
  DFFRX1 \clk_div_reg[10]  ( .D(N249), .CK(n6), .RN(n11), .Q(clk_div[10]) );
  DFFRX1 \clk_div_reg[11]  ( .D(N250), .CK(n6), .RN(n11), .Q(clk_div[11]) );
  DFFRX1 \clk_div_reg[12]  ( .D(N251), .CK(n6), .RN(n11), .Q(clk_div[12]) );
  DFFRX1 \clk_div_reg[1]  ( .D(N240), .CK(n9), .RN(reset_n), .Q(clk_div[1]) );
  DFFRX1 \i_idle_reg[0]  ( .D(n144), .CK(n4), .RN(n2), .Q(i_idle[0]) );
  DFFRX2 \state_reg[0]  ( .D(n146), .CK(n4), .RN(n2), .Q(state[0]), .QN(n8) );
  DFFRXL \i_idle_reg[1]  ( .D(n145), .CK(n4), .RN(n2), .Q(i_idle[1]) );
  DFFRX2 \decoderin1_reg[3]  ( .D(n138), .CK(n4), .RN(n2), .Q(decoderin1[3]), 
        .QN(n12) );
  DFFRX2 \decoderin1_reg[1]  ( .D(n140), .CK(n4), .RN(n2), .Q(decoderin1[1]), 
        .QN(n16) );
  DFFRX2 \decoderin1_reg[2]  ( .D(n139), .CK(n4), .RN(n2), .Q(decoderin1[2]), 
        .QN(n14) );
  DFFRX1 \clk_div_reg[13]  ( .D(N252), .CK(n6), .RN(n11), .Q(clk_div[13]) );
  DFFSX2 \decoderin1_reg[4]  ( .D(n137), .CK(n4), .SN(n2), .Q(decoderin1[4]), 
        .QN(n10) );
  DFFSX2 \decoderin1_reg[0]  ( .D(n141), .CK(n5), .SN(n2), .Q(decoderin1[0]), 
        .QN(n17) );
  NAND4X1 U3 ( .A(i_hex[3]), .B(i_hex[2]), .C(i_hex[1]), .D(i_hex[0]), .Y(n120) );
  OAI211X1 U4 ( .A0(n8), .A1(n120), .B0(n135), .C0(n7), .Y(n134) );
  AOI221XL U5 ( .A0(desOut[37]), .A1(n81), .B0(desOut[33]), .B1(n82), .C0(n123), .Y(n117) );
  AOI221XL U6 ( .A0(desOut[55]), .A1(n77), .B0(desOut[51]), .B1(n78), .C0(n100), .Y(n99) );
  AOI221XL U7 ( .A0(desOut[39]), .A1(n81), .B0(desOut[35]), .B1(n82), .C0(n101), .Y(n98) );
  AOI221XL U8 ( .A0(desOut[54]), .A1(n77), .B0(desOut[50]), .B1(n78), .C0(n109), .Y(n108) );
  AOI221XL U9 ( .A0(desOut[38]), .A1(n81), .B0(desOut[34]), .B1(n82), .C0(n110), .Y(n107) );
  AOI221XL U10 ( .A0(desOut[56]), .A1(n77), .B0(desOut[52]), .B1(n78), .C0(n79), .Y(n76) );
  AOI221XL U11 ( .A0(desOut[40]), .A1(n81), .B0(desOut[36]), .B1(n82), .C0(n83), .Y(n75) );
  OAI222X1 U12 ( .A0(n17), .A1(n71), .B0(n114), .B1(n113), .C0(n27), .C1(n7), 
        .Y(n141) );
  AOI221XL U13 ( .A0(desOut[21]), .A1(n86), .B0(desOut[17]), .B1(n87), .C0(
        n125), .Y(n116) );
  CLKBUFX3 U14 ( .A(clk_div[13]), .Y(n5) );
  CLKBUFX3 U15 ( .A(n90), .Y(n1) );
  NOR3X4 U16 ( .A(n18), .B(i_hex[1]), .C(n124), .Y(n81) );
  NAND2X4 U17 ( .A(i_hex[0]), .B(n21), .Y(n124) );
  NOR4X4 U18 ( .A(i_hex[0]), .B(i_hex[1]), .C(i_hex[2]), .D(i_hex[3]), .Y(n91)
         );
  INVX4 U19 ( .A(n150), .Y(n2) );
  INVX4 U20 ( .A(n150), .Y(n157) );
  NAND2X1 U21 ( .A(desEnable), .B(reset_n), .Y(n150) );
  CLKINVX1 U22 ( .A(n120), .Y(n19) );
  CLKINVX1 U25 ( .A(n126), .Y(n15) );
  NAND2X1 U26 ( .A(n36), .B(n37), .Y(n32) );
  CLKINVX1 U29 ( .A(n39), .Y(n154) );
  CLKINVX1 U30 ( .A(n134), .Y(n20) );
  CLKINVX1 U31 ( .A(n36), .Y(n156) );
  AND2X2 U32 ( .A(n122), .B(n121), .Y(n78) );
  CLKINVX1 U33 ( .A(n62), .Y(n151) );
  CLKINVX1 U34 ( .A(n54), .Y(n152) );
  CLKINVX1 U35 ( .A(n133), .Y(n24) );
  CLKINVX1 U36 ( .A(n63), .Y(n153) );
  CLKINVX1 U37 ( .A(n113), .Y(n29) );
  NAND3X1 U38 ( .A(i_idle[0]), .B(n8), .C(i_idle[1]), .Y(n135) );
  AOI31X1 U39 ( .A0(n35), .A1(n28), .A2(n30), .B0(n39), .Y(n44) );
  NAND3X1 U40 ( .A(decoderin1[4]), .B(n16), .C(n151), .Y(n57) );
  NOR3X1 U41 ( .A(n16), .B(decoderin1[2]), .C(n12), .Y(n65) );
  CLKBUFX3 U42 ( .A(clk_div[13]), .Y(n4) );
  NAND4X1 U43 ( .A(decoderin1[2]), .B(decoderin1[1]), .C(decoderin1[0]), .D(
        n10), .Y(n51) );
  XOR2X1 U44 ( .A(n23), .B(n129), .Y(n149) );
  XNOR2X1 U45 ( .A(i_idle[1]), .B(n132), .Y(n145) );
  NAND2X1 U46 ( .A(n24), .B(i_idle[0]), .Y(n132) );
  XOR2X1 U47 ( .A(i_idle[0]), .B(n24), .Y(n144) );
  NAND3X1 U48 ( .A(n31), .B(n25), .C(decoderin2[2]), .Y(n41) );
  NAND3X1 U49 ( .A(i_hex[2]), .B(i_hex[0]), .C(n127), .Y(n126) );
  NAND3X1 U50 ( .A(n16), .B(n14), .C(n55), .Y(n60) );
  OAI22X1 U51 ( .A0(n126), .A1(n129), .B0(n136), .B1(n18), .Y(n148) );
  NOR2X1 U53 ( .A(n120), .B(n130), .Y(n136) );
  OAI22XL U54 ( .A0(n8), .A1(n134), .B0(n20), .B1(n133), .Y(n146) );
  NOR2X1 U57 ( .A(n129), .B(n23), .Y(n131) );
  OAI2BB2XL U58 ( .B0(n16), .B1(n71), .A0N(n29), .A1N(n104), .Y(n140) );
  NAND4X1 U59 ( .A(n105), .B(n106), .C(n107), .D(n108), .Y(n104) );
  AOI221XL U60 ( .A0(desOut[6]), .A1(n90), .B0(desOut[2]), .B1(n91), .C0(n112), 
        .Y(n105) );
  AOI221XL U61 ( .A0(desOut[22]), .A1(n86), .B0(desOut[18]), .B1(n87), .C0(
        n111), .Y(n106) );
  OAI2BB2XL U62 ( .B0(n14), .B1(n71), .A0N(n29), .A1N(n95), .Y(n139) );
  NAND4X1 U63 ( .A(n96), .B(n97), .C(n98), .D(n99), .Y(n95) );
  AOI221XL U64 ( .A0(desOut[7]), .A1(n90), .B0(desOut[3]), .B1(n91), .C0(n103), 
        .Y(n96) );
  AOI221XL U65 ( .A0(desOut[23]), .A1(n86), .B0(desOut[19]), .B1(n87), .C0(
        n102), .Y(n97) );
  OAI2BB2XL U66 ( .B0(n12), .B1(n71), .A0N(n29), .A1N(n72), .Y(n138) );
  NAND4X1 U67 ( .A(n73), .B(n74), .C(n75), .D(n76), .Y(n72) );
  AOI221XL U68 ( .A0(desOut[8]), .A1(n1), .B0(desOut[4]), .B1(n91), .C0(n92), 
        .Y(n73) );
  AOI221XL U69 ( .A0(desOut[24]), .A1(n86), .B0(desOut[20]), .B1(n87), .C0(n88), .Y(n74) );
  NAND2X1 U70 ( .A(n14), .B(n12), .Y(n62) );
  OAI21XL U71 ( .A0(n10), .A1(n71), .B0(state[0]), .Y(n137) );
  NAND2X1 U72 ( .A(n8), .B(n7), .Y(n133) );
  NAND2X1 U73 ( .A(decoderin1[1]), .B(n17), .Y(n63) );
  NAND2X1 U74 ( .A(n131), .B(i_hex[1]), .Y(n130) );
  NAND2X1 U75 ( .A(state[0]), .B(n71), .Y(n113) );
  OAI211X1 U76 ( .A0(n37), .A1(n45), .B0(n25), .C0(n46), .Y(segout2[2]) );
  NAND2X1 U77 ( .A(n31), .B(n26), .Y(n45) );
  OAI211X1 U78 ( .A0(decoderin2[1]), .A1(n31), .B0(decoderin2[2]), .C0(
        decoderin2[3]), .Y(n46) );
  OAI211X1 U79 ( .A0(decoderin2[1]), .A1(n41), .B0(n50), .C0(n44), .Y(
        segout2[0]) );
  NAND3X1 U80 ( .A(n32), .B(n25), .C(decoderin2[3]), .Y(n50) );
  OAI211X1 U81 ( .A0(n41), .A1(n42), .B0(n43), .C0(n44), .Y(segout2[3]) );
  NAND2X1 U82 ( .A(n30), .B(n26), .Y(n42) );
  NAND4X1 U83 ( .A(decoderin2[0]), .B(decoderin2[2]), .C(decoderin2[1]), .D(
        n25), .Y(n43) );
  OAI211X1 U84 ( .A0(decoderin1[4]), .A1(n69), .B0(n60), .C0(n53), .Y(
        segout1[0]) );
  NOR2X1 U85 ( .A(n61), .B(n65), .Y(n69) );
  OAI211X1 U86 ( .A0(n62), .A1(n63), .B0(n64), .C0(n10), .Y(segout1[2]) );
  OAI211X1 U87 ( .A0(decoderin1[1]), .A1(n17), .B0(decoderin1[2]), .C0(
        decoderin1[3]), .Y(n64) );
  CLKINVX1 U88 ( .A(n70), .Y(n53) );
  OAI31X1 U89 ( .A0(n12), .A1(decoderin1[4]), .A2(n54), .B0(n57), .Y(n70) );
  NAND4BX1 U90 ( .AN(n65), .B(n10), .C(n66), .D(n67), .Y(segout1[1]) );
  NAND3X1 U91 ( .A(decoderin1[2]), .B(n12), .C(n153), .Y(n66) );
  AOI22X1 U92 ( .A0(decoderin1[3]), .A1(n68), .B0(n55), .B1(n152), .Y(n67) );
  AO21X1 U94 ( .A0(decoderin1[0]), .A1(decoderin1[1]), .B0(n61), .Y(n68) );
  NAND4X1 U96 ( .A(n59), .B(n51), .C(n60), .D(n57), .Y(segout1[3]) );
  NAND3X1 U97 ( .A(n12), .B(n10), .C(n61), .Y(n59) );
  NOR2X1 U102 ( .A(n8), .B(n20), .Y(n147) );
  NOR3X1 U103 ( .A(n32), .B(decoderin2[3]), .C(n33), .Y(segout2[6]) );
  AOI2BB2X1 U104 ( .B0(decoderin2[0]), .B1(n25), .A0N(decoderin2[0]), .A1N(
        decoderin2[1]), .Y(n33) );
  OAI21XL U109 ( .A0(decoderin1[3]), .A1(n51), .B0(n52), .Y(segout1[6]) );
  OAI211X1 U110 ( .A0(n17), .A1(n10), .B0(n16), .C0(n151), .Y(n52) );
  OAI21XL U113 ( .A0(decoderin1[4]), .A1(n56), .B0(n57), .Y(segout1[4]) );
  AOI21XL U116 ( .A0(n58), .A1(n16), .B0(n55), .Y(n56) );
  OAI22X1 U117 ( .A0(decoderin1[3]), .A1(n14), .B0(decoderin1[2]), .B1(n17), 
        .Y(n58) );
  OAI21XL U118 ( .A0(decoderin2[4]), .A1(n38), .B0(n154), .Y(segout2[4]) );
  AOI21X1 U119 ( .A0(n40), .A1(n30), .B0(n35), .Y(n38) );
  OAI22X1 U120 ( .A0(decoderin2[3]), .A1(n28), .B0(decoderin2[2]), .B1(n31), 
        .Y(n40) );
  OAI21XL U121 ( .A0(decoderin2[4]), .A1(n34), .B0(n154), .Y(segout2[5]) );
  AOI222XL U122 ( .A0(decoderin2[3]), .A1(n156), .B0(n155), .B1(n31), .C0(n35), 
        .C1(n36), .Y(n34) );
  CLKINVX1 U123 ( .A(n37), .Y(n155) );
  NAND3X1 U124 ( .A(n47), .B(n25), .C(n48), .Y(segout2[1]) );
  AOI22XL U125 ( .A0(n156), .A1(n35), .B0(decoderin2[3]), .B1(n49), .Y(n48) );
  NAND4X1 U126 ( .A(decoderin2[2]), .B(decoderin2[1]), .C(n31), .D(n26), .Y(
        n47) );
  OAI221X1 U127 ( .A0(decoderin2[0]), .A1(n36), .B0(n30), .B1(n31), .C0(n37), 
        .Y(n49) );
  BUFX4 U128 ( .A(reset_n), .Y(n11) );
  AO22X1 U129 ( .A0(desOut[58]), .A1(n80), .B0(desOut[62]), .B1(n19), .Y(n109)
         );
  AO22X1 U130 ( .A0(desOut[59]), .A1(n80), .B0(desOut[63]), .B1(n19), .Y(n100)
         );
  AO22X1 U131 ( .A0(desOut[60]), .A1(n80), .B0(desOut[64]), .B1(n19), .Y(n79)
         );
  AO22X1 U132 ( .A0(desOut[42]), .A1(n84), .B0(desOut[46]), .B1(n85), .Y(n110)
         );
  AO22XL U134 ( .A0(desOut[43]), .A1(n84), .B0(desOut[47]), .B1(n85), .Y(n101)
         );
  AO22XL U136 ( .A0(desOut[44]), .A1(n84), .B0(desOut[48]), .B1(n85), .Y(n83)
         );
  AOI221XL U137 ( .A0(desOut[53]), .A1(n77), .B0(desOut[49]), .B1(n78), .C0(
        n119), .Y(n118) );
  AO22X1 U138 ( .A0(desOut[57]), .A1(n80), .B0(desOut[61]), .B1(n19), .Y(n119)
         );
  AND4X1 U139 ( .A(n115), .B(n116), .C(n117), .D(n118), .Y(n114) );
  INVXL U140 ( .A(n71), .Y(n27) );
  AOI221XL U141 ( .A0(desOut[5]), .A1(n1), .B0(desOut[1]), .B1(n91), .C0(n128), 
        .Y(n115) );
  AO22XL U142 ( .A0(desOut[41]), .A1(n84), .B0(desOut[45]), .B1(n85), .Y(n123)
         );
  AO22X1 U143 ( .A0(desOut[25]), .A1(n89), .B0(desOut[29]), .B1(n15), .Y(n125)
         );
  AO22X1 U144 ( .A0(desOut[9]), .A1(n93), .B0(desOut[13]), .B1(n94), .Y(n128)
         );
  AO22X1 U145 ( .A0(desOut[26]), .A1(n89), .B0(desOut[30]), .B1(n15), .Y(n111)
         );
  AO22X1 U146 ( .A0(desOut[10]), .A1(n93), .B0(desOut[14]), .B1(n94), .Y(n112)
         );
  AO22X1 U147 ( .A0(desOut[27]), .A1(n89), .B0(desOut[31]), .B1(n15), .Y(n102)
         );
  AO22X1 U148 ( .A0(desOut[11]), .A1(n93), .B0(desOut[15]), .B1(n94), .Y(n103)
         );
  AO22X1 U149 ( .A0(desOut[28]), .A1(n89), .B0(desOut[32]), .B1(n15), .Y(n88)
         );
  AO22X1 U150 ( .A0(desOut[12]), .A1(n93), .B0(desOut[16]), .B1(n94), .Y(n92)
         );
  OAI21XL U151 ( .A0(n3), .A1(decoderin1[4]), .B0(n53), .Y(segout1[5]) );
  AOI22X1 U152 ( .A0(n14), .A1(n153), .B0(n54), .B1(n55), .Y(n3) );
  OAI32X1 U153 ( .A0(n129), .A1(n22), .A2(n124), .B0(n13), .B1(n21), .Y(n142)
         );
  CLKINVX1 U154 ( .A(n130), .Y(n13) );
  OAI32X1 U155 ( .A0(n129), .A1(i_hex[1]), .A2(n23), .B0(n131), .B1(n22), .Y(
        n143) );
  CLKBUFX3 U156 ( .A(clk), .Y(n6) );
  CLKBUFX3 U157 ( .A(clk), .Y(n9) );
endmodule


module des2_top ( dip1, dip2, dip3, dip4, dip5, dip6, dip7, dip8, dip9, 
        reset_n, clk, segout1, segout2 );
  output [6:0] segout1;
  output [6:0] segout2;
  input dip1, dip2, dip3, dip4, dip5, dip6, dip7, dip8, dip9, reset_n, clk;
  wire   decrypt, desEnable;
  wire   [3:1] key1sel;
  wire   [3:1] key2sel;
  wire   [63:0] desIn;
  wire   [55:0] key1;
  wire   [55:0] key2;
  wire   [63:0] desOut;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103;

  dip_driver DIP ( .dip1(dip1), .dip2(dip2), .dip3(dip3), .dip4(dip4), .dip5(
        dip5), .dip6(dip6), .dip7(dip7), .dip8(dip8), .dip9(dip9), .reset_n(
        reset_n), .key1sel(key1sel), .key2sel(key2sel), .decrypt(decrypt), 
        .desEnable(desEnable), .desIn(desIn) );
  keybox KBX ( .key1sel(key1sel), .key2sel(key2sel), .key1({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, key1[47:44], 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51}), .key2({
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, key2[47:44], 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103}) );
  des2 DES ( .desIn(desIn), .key1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, key1[47:44], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .key2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, key2[47:44], 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .decrypt(decrypt), 
        .desEnable(desEnable), .reset_n(reset_n), .clk(clk), .desOut(desOut)
         );
  seg_decoder SEG ( .desOut(desOut), .desEnable(desEnable), .reset_n(reset_n), 
        .clk(clk), .segout1(segout1), .segout2(segout2) );
endmodule

